magic
tech sky130A
timestamp 1765331190
<< error_s >>
rect -110 295 85 440
rect -340 140 85 295
rect -320 5 -285 55
rect -270 5 -235 55
rect -205 5 -170 55
rect -155 5 -120 55
rect -90 5 -45 55
rect -30 5 15 55
rect 30 5 65 55
rect -90 -90 -75 5
rect 50 -90 65 5
rect -90 -140 -45 -90
rect -30 -140 -5 -90
rect 10 -140 65 -90
<< nwell >>
rect -110 140 85 440
<< nmos >>
rect -45 5 -30 55
rect 15 5 30 55
rect -45 -140 -30 -90
rect -5 -140 10 -90
<< pmos >>
rect -45 370 -30 420
rect 15 370 30 420
rect -45 225 -30 275
rect 15 225 30 275
<< ndiff >>
rect -90 5 -45 55
rect -30 5 15 55
rect 30 5 65 55
rect -90 -90 -75 5
rect 50 -90 65 5
rect -90 -105 -45 -90
rect -90 -125 -85 -105
rect -65 -125 -45 -105
rect -90 -140 -45 -125
rect -30 -140 -5 -90
rect 10 -100 65 -90
rect 10 -120 35 -100
rect 55 -120 65 -100
rect 10 -140 65 -120
<< pdiff >>
rect -90 405 -45 420
rect -90 385 -85 405
rect -65 385 -45 405
rect -90 370 -45 385
rect -30 370 15 420
rect 30 370 65 420
rect -90 275 -75 370
rect 50 275 65 370
rect -90 225 -45 275
rect -30 225 15 275
rect 30 260 65 275
rect 30 240 40 260
rect 60 240 65 260
rect 30 225 65 240
<< ndiffc >>
rect -85 -125 -65 -105
rect 35 -120 55 -100
<< pdiffc >>
rect -85 385 -65 405
rect 40 240 60 260
<< poly >>
rect -45 420 -30 435
rect 15 420 30 435
rect -45 355 -30 370
rect 15 355 30 370
rect -55 345 -25 355
rect -55 325 -50 345
rect -30 325 -25 345
rect -55 315 -25 325
rect 0 345 30 355
rect 0 325 5 345
rect 25 325 30 345
rect 0 315 30 325
rect -45 275 -30 290
rect 15 275 30 290
rect -45 200 -30 225
rect 15 210 30 225
rect -170 185 -30 200
rect -45 140 -30 185
rect -5 200 30 210
rect -5 180 0 200
rect 20 180 30 200
rect -5 170 30 180
rect -45 125 30 140
rect -90 95 -60 105
rect -90 75 -85 95
rect -65 80 -60 95
rect -65 75 -30 80
rect -90 65 -30 75
rect -45 55 -30 65
rect 15 55 30 125
rect -45 -10 -30 5
rect 15 -10 30 5
rect -60 -45 -30 -35
rect -60 -65 -55 -45
rect -35 -65 -30 -45
rect -60 -75 -30 -65
rect -45 -90 -30 -75
rect -5 -45 30 -35
rect -5 -65 0 -45
rect 20 -65 30 -45
rect -5 -75 30 -65
rect -5 -90 10 -75
rect -45 -155 -30 -140
rect -5 -155 10 -140
<< polycont >>
rect -50 325 -30 345
rect 5 325 25 345
rect 0 180 20 200
rect -85 75 -65 95
rect -55 -65 -35 -45
rect 0 -65 20 -45
<< locali >>
rect -90 405 -60 420
rect -90 395 -85 405
rect -125 385 -85 395
rect -65 385 -60 405
rect -125 375 -60 385
rect -125 310 -105 375
rect -55 345 -25 355
rect -55 335 -50 345
rect -310 290 -105 310
rect -85 325 -50 335
rect -30 325 -25 345
rect -85 315 -25 325
rect -5 345 30 355
rect -5 325 5 345
rect 25 325 30 345
rect -5 315 30 325
rect -310 275 -290 290
rect -205 275 -175 290
rect -320 180 -185 200
rect -205 120 -185 180
rect -305 100 -285 120
rect -85 105 -65 315
rect -5 250 15 315
rect -45 230 15 250
rect 35 260 65 275
rect 35 240 40 260
rect 60 240 65 260
rect -45 150 -25 230
rect 35 225 65 240
rect -5 200 25 210
rect -5 180 0 200
rect 20 180 25 200
rect -5 170 25 180
rect -45 130 -15 150
rect -90 100 -60 105
rect -320 95 -60 100
rect -320 80 -85 95
rect -90 75 -85 80
rect -65 75 -60 95
rect -90 65 -60 75
rect -35 45 -15 130
rect -120 25 -15 45
rect -35 5 -15 25
rect -310 -10 -290 5
rect -205 -10 -175 5
rect -310 -30 -80 -10
rect -100 -95 -80 -30
rect -45 -15 -15 5
rect -45 -35 -25 -15
rect 5 -35 25 170
rect -60 -45 -25 -35
rect -60 -65 -55 -45
rect -35 -65 -25 -45
rect -60 -75 -25 -65
rect -5 -45 25 -35
rect -5 -65 0 -45
rect 20 -65 25 -45
rect -5 -75 25 -65
rect 45 -95 65 225
rect -100 -105 -60 -95
rect -100 -125 -85 -105
rect -65 -125 -60 -105
rect 25 -100 65 -95
rect 25 -120 35 -100
rect 55 -120 65 -100
rect 25 -125 65 -120
rect -100 -140 -60 -125
<< viali >>
rect 0 -65 20 -45
<< metal1 >>
rect -255 -10 -235 10
rect -255 -30 25 -10
rect -5 -45 25 -30
rect -5 -65 0 -45
rect 20 -65 25 -45
rect -5 -75 25 -65
use inv  inv_0
timestamp 1765330272
transform 1 0 -185 0 1 0
box -40 -10 85 295
use inv  inv_1
timestamp 1765330272
transform 1 0 -300 0 1 0
box -40 -10 85 295
<< end >>
