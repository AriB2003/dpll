magic
tech sky130A
timestamp 1765141373
<< nwell >>
rect -25 300 65 400
rect -40 295 65 300
rect -40 140 85 295
<< nmos >>
rect 15 5 30 55
<< pmos >>
rect 15 225 30 275
<< ndiff >>
rect -20 40 15 55
rect -20 20 -15 40
rect 5 20 15 40
rect -20 5 15 20
rect 30 40 65 55
rect 30 20 40 40
rect 60 20 65 40
rect 30 5 65 20
<< pdiff >>
rect -20 260 15 275
rect -20 240 -15 260
rect 5 240 15 260
rect -20 225 15 240
rect 30 260 65 275
rect 30 240 40 260
rect 60 240 65 260
rect 30 225 65 240
<< ndiffc >>
rect -15 20 5 40
rect 40 20 60 40
<< pdiffc >>
rect -15 240 5 260
rect 40 240 60 260
<< psubdiff >>
rect 0 -40 50 -25
rect 0 -65 15 -40
rect 35 -65 50 -40
rect 0 -80 50 -65
<< nsubdiff >>
rect -5 365 45 380
rect -5 340 10 365
rect 30 340 45 365
rect -5 325 45 340
<< psubdiffcont >>
rect 15 -65 35 -40
<< nsubdiffcont >>
rect 10 340 30 365
<< poly >>
rect 15 275 30 290
rect 15 160 30 225
rect -15 150 30 160
rect -15 130 -10 150
rect 10 130 30 150
rect -15 120 30 130
rect 15 55 30 120
rect 15 -10 30 5
<< polycont >>
rect -10 130 10 150
<< locali >>
rect 5 365 35 375
rect 5 340 10 365
rect 30 340 35 365
rect 5 330 35 340
rect -20 260 10 275
rect -20 240 -15 260
rect 5 240 10 260
rect -20 225 10 240
rect 35 260 65 275
rect 35 240 40 260
rect 60 240 65 260
rect 35 225 65 240
rect -15 150 15 160
rect -20 130 -10 150
rect 10 130 15 150
rect -15 120 15 130
rect 35 150 65 160
rect 35 130 40 150
rect 60 130 65 150
rect 35 120 65 130
rect -20 40 10 55
rect -20 20 -15 40
rect 5 20 10 40
rect -20 5 10 20
rect 35 40 65 55
rect 35 20 40 40
rect 60 20 65 40
rect 35 5 65 20
rect 10 -40 40 -30
rect 10 -65 15 -40
rect 35 -65 40 -40
rect 10 -75 40 -65
<< viali >>
rect 40 240 60 260
rect 40 130 60 150
rect 40 20 60 40
<< metal1 >>
rect 35 260 65 275
rect 35 240 40 260
rect 60 240 65 260
rect 35 150 65 240
rect 35 130 40 150
rect 60 130 65 150
rect 35 40 65 130
rect 35 20 40 40
rect 60 20 65 40
rect 35 5 65 20
<< end >>
