magic
tech sky130A
timestamp 1765329033
<< nwell >>
rect 2750 505 2895 605
rect 120 400 2895 455
rect -25 310 2895 400
rect -140 300 2895 310
rect -1000 290 2895 300
rect -1000 160 70 290
rect 270 230 300 290
rect 470 230 500 290
rect 670 230 700 290
rect 870 230 900 290
rect 1070 230 1100 290
rect 1270 230 1300 290
rect 1470 230 1500 290
rect 1670 230 1700 290
rect 1870 230 1900 290
rect 2070 230 2100 290
rect 2270 230 2300 290
rect 2470 230 2500 290
rect 2670 230 2700 290
rect 2790 230 2820 290
rect -1000 140 95 160
<< nmos >>
rect -945 5 -895 55
rect -855 5 -805 55
rect -765 5 -715 55
rect -675 5 -625 55
rect -585 5 -535 55
rect -495 5 -445 55
rect -405 5 -355 55
rect -315 5 -265 55
rect -225 5 -175 55
rect -135 5 -85 55
rect 15 5 65 55
<< pmos >>
rect -945 225 -895 275
rect -855 225 -805 275
rect -765 225 -715 275
rect -675 225 -625 275
rect -585 225 -535 275
rect -495 225 -445 275
rect -405 225 -355 275
rect -315 225 -265 275
rect -225 225 -175 275
rect -135 225 -85 275
rect 15 225 65 275
<< ndiff >>
rect -980 40 -945 55
rect -980 20 -975 40
rect -955 20 -945 40
rect -980 5 -945 20
rect -895 40 -855 55
rect -895 20 -885 40
rect -865 20 -855 40
rect -895 5 -855 20
rect -805 40 -765 55
rect -805 20 -795 40
rect -775 20 -765 40
rect -805 5 -765 20
rect -715 40 -675 55
rect -715 20 -705 40
rect -685 20 -675 40
rect -715 5 -675 20
rect -625 40 -585 55
rect -625 20 -615 40
rect -595 20 -585 40
rect -625 5 -585 20
rect -535 40 -495 55
rect -535 20 -525 40
rect -505 20 -495 40
rect -535 5 -495 20
rect -445 40 -405 55
rect -445 20 -435 40
rect -415 20 -405 40
rect -445 5 -405 20
rect -355 40 -315 55
rect -355 20 -345 40
rect -325 20 -315 40
rect -355 5 -315 20
rect -265 40 -225 55
rect -265 20 -255 40
rect -235 20 -225 40
rect -265 5 -225 20
rect -175 40 -135 55
rect -175 20 -165 40
rect -145 20 -135 40
rect -175 5 -135 20
rect -85 40 -50 55
rect -85 20 -75 40
rect -55 20 -50 40
rect -85 5 -50 20
rect -20 40 15 55
rect -20 20 -15 40
rect 5 20 15 40
rect -20 5 15 20
rect 65 5 70 55
<< pdiff >>
rect -980 260 -945 275
rect -980 240 -975 260
rect -955 240 -945 260
rect -980 225 -945 240
rect -895 260 -855 275
rect -895 240 -885 260
rect -865 240 -855 260
rect -895 225 -855 240
rect -805 260 -765 275
rect -805 240 -795 260
rect -775 240 -765 260
rect -805 225 -765 240
rect -715 260 -675 275
rect -715 240 -705 260
rect -685 240 -675 260
rect -715 225 -675 240
rect -625 260 -585 275
rect -625 240 -615 260
rect -595 240 -585 260
rect -625 225 -585 240
rect -535 260 -495 275
rect -535 240 -525 260
rect -505 240 -495 260
rect -535 225 -495 240
rect -445 260 -405 275
rect -445 240 -435 260
rect -415 240 -405 260
rect -445 225 -405 240
rect -355 260 -315 275
rect -355 240 -345 260
rect -325 240 -315 260
rect -355 225 -315 240
rect -265 260 -225 275
rect -265 240 -255 260
rect -235 240 -225 260
rect -265 225 -225 240
rect -175 260 -135 275
rect -175 240 -165 260
rect -145 240 -135 260
rect -175 225 -135 240
rect -85 260 -50 275
rect -85 240 -75 260
rect -55 240 -50 260
rect -85 225 -50 240
rect -20 260 15 275
rect -20 240 -15 260
rect 5 240 15 260
rect -20 225 15 240
rect 65 225 70 275
<< ndiffc >>
rect -975 20 -955 40
rect -885 20 -865 40
rect -795 20 -775 40
rect -705 20 -685 40
rect -615 20 -595 40
rect -525 20 -505 40
rect -435 20 -415 40
rect -345 20 -325 40
rect -255 20 -235 40
rect -165 20 -145 40
rect -75 20 -55 40
rect -15 20 5 40
<< pdiffc >>
rect -975 240 -955 260
rect -885 240 -865 260
rect -795 240 -775 260
rect -705 240 -685 260
rect -615 240 -595 260
rect -525 240 -505 260
rect -435 240 -415 260
rect -345 240 -325 260
rect -255 240 -235 260
rect -165 240 -145 260
rect -75 240 -55 260
rect -15 240 5 260
<< psubdiff >>
rect 0 -40 50 -25
rect 0 -65 15 -40
rect 35 -65 50 -40
rect 0 -80 50 -65
<< nsubdiff >>
rect -5 365 45 380
rect -5 340 10 365
rect 30 340 45 365
rect -5 325 45 340
<< psubdiffcont >>
rect 15 -65 35 -40
<< nsubdiffcont >>
rect 10 340 30 365
<< poly >>
rect -945 275 -895 290
rect -855 275 -805 290
rect -765 275 -715 290
rect -675 275 -625 290
rect -585 275 -535 290
rect -495 275 -445 290
rect -405 275 -355 290
rect -315 275 -265 290
rect -225 275 -175 290
rect -135 275 -85 290
rect 15 275 65 290
rect -945 210 -895 225
rect -855 210 -805 225
rect -765 210 -715 225
rect -675 210 -625 225
rect -585 210 -535 225
rect -495 210 -445 225
rect -405 210 -355 225
rect -315 210 -265 225
rect -225 210 -175 225
rect -135 210 -85 225
rect 15 210 65 225
rect -935 200 -905 210
rect -935 180 -930 200
rect -910 180 -905 200
rect -935 170 -905 180
rect -845 200 -815 210
rect -845 180 -840 200
rect -820 180 -815 200
rect -845 170 -815 180
rect -755 200 -725 210
rect -755 180 -750 200
rect -730 180 -725 200
rect -755 170 -725 180
rect -665 200 -635 210
rect -665 180 -660 200
rect -640 180 -635 200
rect -665 170 -635 180
rect -575 200 -545 210
rect -575 180 -570 200
rect -550 180 -545 200
rect -575 170 -545 180
rect -485 200 -455 210
rect -485 180 -480 200
rect -460 180 -455 200
rect -485 170 -455 180
rect -395 200 -365 210
rect -395 180 -390 200
rect -370 180 -365 200
rect -395 170 -365 180
rect -305 200 -275 210
rect -305 180 -300 200
rect -280 180 -275 200
rect -305 170 -275 180
rect -215 200 -185 210
rect -215 180 -210 200
rect -190 180 -185 200
rect -215 170 -185 180
rect -125 200 -95 210
rect -125 180 -120 200
rect -100 180 -95 200
rect -125 170 -95 180
rect 20 200 50 210
rect 20 180 25 200
rect 45 180 50 200
rect 20 170 50 180
rect -935 100 -905 110
rect -935 80 -930 100
rect -910 80 -905 100
rect -935 70 -905 80
rect -845 100 -815 110
rect -845 80 -840 100
rect -820 80 -815 100
rect -845 70 -815 80
rect -755 100 -725 110
rect -755 80 -750 100
rect -730 80 -725 100
rect -755 70 -725 80
rect -665 100 -635 110
rect -665 80 -660 100
rect -640 80 -635 100
rect -665 70 -635 80
rect -575 100 -545 110
rect -575 80 -570 100
rect -550 80 -545 100
rect -575 70 -545 80
rect -485 100 -455 110
rect -485 80 -480 100
rect -460 80 -455 100
rect -485 70 -455 80
rect -395 100 -365 110
rect -395 80 -390 100
rect -370 80 -365 100
rect -395 70 -365 80
rect -305 100 -275 110
rect -305 80 -300 100
rect -280 80 -275 100
rect -305 70 -275 80
rect -215 100 -185 110
rect -215 80 -210 100
rect -190 80 -185 100
rect -215 70 -185 80
rect -125 100 -95 110
rect -125 80 -120 100
rect -100 80 -95 100
rect -125 70 -95 80
rect 20 100 50 110
rect 20 80 25 100
rect 45 80 50 100
rect 20 70 50 80
rect -945 55 -895 70
rect -855 55 -805 70
rect -765 55 -715 70
rect -675 55 -625 70
rect -585 55 -535 70
rect -495 55 -445 70
rect -405 55 -355 70
rect -315 55 -265 70
rect -225 55 -175 70
rect -135 55 -85 70
rect 15 55 65 70
rect -945 -10 -895 5
rect -855 -10 -805 5
rect -765 -10 -715 5
rect -675 -10 -625 5
rect -585 -10 -535 5
rect -495 -10 -445 5
rect -405 -10 -355 5
rect -315 -10 -265 5
rect -225 -10 -175 5
rect -135 -10 -85 5
rect 15 -10 65 5
<< polycont >>
rect -930 180 -910 200
rect -840 180 -820 200
rect -750 180 -730 200
rect -660 180 -640 200
rect -570 180 -550 200
rect -480 180 -460 200
rect -390 180 -370 200
rect -300 180 -280 200
rect -210 180 -190 200
rect -120 180 -100 200
rect 25 180 45 200
rect -930 80 -910 100
rect -840 80 -820 100
rect -750 80 -730 100
rect -660 80 -640 100
rect -570 80 -550 100
rect -480 80 -460 100
rect -390 80 -370 100
rect -300 80 -280 100
rect -210 80 -190 100
rect -120 80 -100 100
rect 25 80 45 100
<< locali >>
rect 5 365 35 375
rect 5 340 10 365
rect 30 340 35 365
rect 5 330 35 340
rect -980 260 -950 275
rect -980 240 -975 260
rect -955 240 -950 260
rect -980 225 -950 240
rect -890 260 -860 275
rect -890 240 -885 260
rect -865 240 -860 260
rect -890 225 -860 240
rect -800 260 -770 275
rect -800 240 -795 260
rect -775 240 -770 260
rect -800 225 -770 240
rect -710 260 -680 275
rect -710 240 -705 260
rect -685 240 -680 260
rect -710 225 -680 240
rect -620 260 -590 275
rect -620 240 -615 260
rect -595 240 -590 260
rect -620 225 -590 240
rect -530 260 -500 275
rect -530 240 -525 260
rect -505 240 -500 260
rect -530 225 -500 240
rect -440 260 -410 275
rect -440 240 -435 260
rect -415 240 -410 260
rect -440 225 -410 240
rect -350 260 -320 275
rect -350 240 -345 260
rect -325 240 -320 260
rect -350 225 -320 240
rect -260 260 -230 275
rect -260 240 -255 260
rect -235 240 -230 260
rect -260 225 -230 240
rect -170 260 -140 275
rect -170 240 -165 260
rect -145 240 -140 260
rect -170 225 -140 240
rect -80 260 -50 275
rect -80 240 -75 260
rect -55 240 -50 260
rect -80 225 -50 240
rect -20 260 10 270
rect -20 240 -15 260
rect 5 240 10 260
rect -20 225 10 240
rect -975 200 -955 225
rect -935 200 -905 210
rect -845 200 -815 210
rect -795 200 -775 225
rect -755 200 -725 210
rect -665 200 -635 210
rect -615 200 -595 225
rect -575 200 -545 210
rect -485 200 -455 210
rect -435 200 -415 225
rect -395 200 -365 210
rect -305 200 -275 210
rect -255 200 -235 225
rect -215 200 -185 210
rect -125 200 -95 210
rect -75 200 -55 225
rect 20 200 50 210
rect -975 180 -930 200
rect -910 180 -840 200
rect -820 180 -750 200
rect -730 180 -660 200
rect -640 180 -570 200
rect -550 180 -480 200
rect -460 180 -390 200
rect -370 180 -300 200
rect -280 180 -210 200
rect -190 180 -120 200
rect -100 180 25 200
rect 45 180 70 200
rect 240 180 275 200
rect 440 180 475 200
rect 640 180 675 200
rect 840 180 875 200
rect 1040 180 1075 200
rect 1240 180 1275 200
rect 1440 180 1475 200
rect 1640 180 1675 200
rect 1840 180 1875 200
rect 2040 180 2075 200
rect 2240 180 2275 200
rect 2440 180 2475 200
rect -975 55 -955 180
rect -935 170 -905 180
rect -845 170 -815 180
rect -935 100 -905 110
rect -845 100 -815 110
rect -935 80 -930 100
rect -910 80 -840 100
rect -820 80 -815 100
rect -935 70 -905 80
rect -845 70 -815 80
rect -795 55 -775 180
rect -755 170 -725 180
rect -665 170 -635 180
rect -755 100 -725 110
rect -665 100 -635 110
rect -755 80 -750 100
rect -730 80 -660 100
rect -640 80 -635 100
rect -755 70 -725 80
rect -665 70 -635 80
rect -615 55 -595 180
rect -575 170 -545 180
rect -485 170 -455 180
rect -575 100 -545 110
rect -485 100 -455 110
rect -575 80 -570 100
rect -550 80 -480 100
rect -460 80 -455 100
rect -575 70 -545 80
rect -485 70 -455 80
rect -435 55 -415 180
rect -395 170 -365 180
rect -305 170 -275 180
rect -395 100 -365 110
rect -305 100 -275 110
rect -395 80 -390 100
rect -370 80 -300 100
rect -280 80 -275 100
rect -395 70 -365 80
rect -305 70 -275 80
rect -255 55 -235 180
rect -215 170 -185 180
rect -125 170 -95 180
rect -215 100 -185 110
rect -125 100 -95 110
rect -215 80 -210 100
rect -190 80 -120 100
rect -100 80 -95 100
rect -215 70 -185 80
rect -125 70 -95 80
rect -75 55 -55 180
rect 20 170 50 180
rect 65 150 95 160
rect 65 130 70 150
rect 90 130 95 150
rect 240 130 275 150
rect 440 130 475 150
rect 640 130 675 150
rect 840 130 875 150
rect 1040 130 1075 150
rect 1240 130 1275 150
rect 1440 130 1475 150
rect 1640 130 1675 150
rect 1840 130 1875 150
rect 2040 130 2075 150
rect 2240 130 2275 150
rect 2440 130 2475 150
rect 2635 130 2670 150
rect 2755 130 2790 150
rect 65 120 95 130
rect 20 100 50 110
rect 20 80 25 100
rect 45 80 70 100
rect 240 80 275 100
rect 440 80 475 100
rect 640 80 675 100
rect 840 80 875 100
rect 1040 80 1075 100
rect 1240 80 1275 100
rect 1440 80 1475 100
rect 1640 80 1675 100
rect 1840 80 1875 100
rect 2040 80 2075 100
rect 2240 80 2275 100
rect 2440 80 2475 100
rect 20 70 50 80
rect -980 40 -950 55
rect -980 20 -975 40
rect -955 20 -950 40
rect -980 10 -950 20
rect -890 40 -860 55
rect -890 20 -885 40
rect -865 20 -860 40
rect -890 10 -860 20
rect -800 40 -770 55
rect -800 20 -795 40
rect -775 20 -770 40
rect -800 10 -770 20
rect -710 40 -680 55
rect -710 20 -705 40
rect -685 20 -680 40
rect -710 10 -680 20
rect -620 40 -590 55
rect -620 20 -615 40
rect -595 20 -590 40
rect -620 10 -590 20
rect -530 40 -500 55
rect -530 20 -525 40
rect -505 20 -500 40
rect -530 10 -500 20
rect -440 40 -410 55
rect -440 20 -435 40
rect -415 20 -410 40
rect -440 10 -410 20
rect -350 40 -320 55
rect -350 20 -345 40
rect -325 20 -320 40
rect -350 10 -320 20
rect -260 40 -230 55
rect -260 20 -255 40
rect -235 20 -230 40
rect -260 10 -230 20
rect -170 40 -140 55
rect -170 20 -165 40
rect -145 20 -140 40
rect -170 10 -140 20
rect -80 40 -50 55
rect -80 20 -75 40
rect -55 20 -50 40
rect -80 10 -50 20
rect -20 40 10 55
rect -20 20 -15 40
rect 5 20 10 40
rect -20 10 10 20
rect 10 -40 40 -30
rect 10 -65 15 -40
rect 35 -65 40 -40
rect 10 -75 40 -65
<< viali >>
rect -885 240 -865 260
rect -705 240 -685 260
rect -525 240 -505 260
rect -345 240 -325 260
rect -165 240 -145 260
rect -15 240 5 260
rect 75 240 95 260
rect 275 240 295 260
rect 475 240 495 260
rect 675 240 695 260
rect 875 240 895 260
rect 1075 240 1095 260
rect 1275 240 1295 260
rect 1475 240 1495 260
rect 1675 240 1695 260
rect 1875 240 1895 260
rect 2075 240 2095 260
rect 2275 240 2295 260
rect 2475 240 2495 260
rect 2675 240 2695 260
rect 2795 240 2815 260
rect -930 80 -910 100
rect -750 80 -730 100
rect -570 80 -550 100
rect -390 80 -370 100
rect -210 80 -190 100
rect 70 130 90 150
rect 25 80 45 100
rect -885 20 -865 40
rect -705 20 -685 40
rect -525 20 -505 40
rect -345 20 -325 40
rect -165 20 -145 40
rect -15 20 5 40
rect 75 20 95 40
rect 275 20 295 40
rect 475 20 495 40
rect 675 20 695 40
rect 875 20 895 40
rect 1075 20 1095 40
rect 1275 20 1295 40
rect 1475 20 1495 40
rect 1675 20 1695 40
rect 1875 20 1895 40
rect 2075 20 2095 40
rect 2275 20 2295 40
rect 2475 20 2495 40
rect 2675 20 2695 40
rect 2795 20 2815 40
<< metal1 >>
rect -170 290 2820 310
rect -890 260 -860 275
rect -710 260 -680 275
rect -530 260 -500 275
rect -350 260 -320 275
rect -170 260 -140 290
rect 70 270 90 290
rect -890 240 -885 260
rect -865 240 -705 260
rect -685 240 -525 260
rect -505 240 -345 260
rect -325 240 -165 260
rect -145 240 -140 260
rect -890 225 -860 240
rect -710 225 -680 240
rect -530 225 -500 240
rect -350 225 -320 240
rect -170 225 -140 240
rect -20 260 10 270
rect -20 240 -15 260
rect 5 240 10 260
rect -20 110 10 240
rect 70 260 100 270
rect 70 240 75 260
rect 95 240 100 260
rect 70 230 100 240
rect 270 260 300 290
rect 270 240 275 260
rect 295 240 300 260
rect 270 230 300 240
rect 470 260 500 290
rect 470 240 475 260
rect 495 240 500 260
rect 470 230 500 240
rect 670 260 700 290
rect 670 240 675 260
rect 695 240 700 260
rect 670 230 700 240
rect 870 260 900 290
rect 870 240 875 260
rect 895 240 900 260
rect 870 230 900 240
rect 1070 260 1100 290
rect 1070 240 1075 260
rect 1095 240 1100 260
rect 1070 230 1100 240
rect 1270 260 1300 290
rect 1270 240 1275 260
rect 1295 240 1300 260
rect 1270 230 1300 240
rect 1470 260 1500 290
rect 1470 240 1475 260
rect 1495 240 1500 260
rect 1470 230 1500 240
rect 1670 260 1700 290
rect 1670 240 1675 260
rect 1695 240 1700 260
rect 1670 230 1700 240
rect 1870 260 1900 290
rect 1870 240 1875 260
rect 1895 240 1900 260
rect 1870 230 1900 240
rect 2070 260 2100 290
rect 2070 240 2075 260
rect 2095 240 2100 260
rect 2070 230 2100 240
rect 2270 260 2300 290
rect 2270 240 2275 260
rect 2295 240 2300 260
rect 2270 230 2300 240
rect 2470 260 2500 290
rect 2470 240 2475 260
rect 2495 240 2500 260
rect 2470 230 2500 240
rect 2670 260 2700 290
rect 2670 240 2675 260
rect 2695 240 2700 260
rect 2670 230 2700 240
rect 2790 260 2820 290
rect 2790 240 2795 260
rect 2815 240 2820 260
rect 2790 230 2820 240
rect 65 155 95 160
rect 65 120 95 125
rect -935 100 -905 110
rect -755 100 -725 110
rect -575 100 -545 110
rect -395 100 -365 110
rect -215 100 -185 110
rect -935 80 -930 100
rect -910 80 -750 100
rect -730 80 -570 100
rect -550 80 -390 100
rect -370 80 -210 100
rect -190 80 -185 100
rect -935 70 -905 80
rect -755 70 -725 80
rect -575 70 -545 80
rect -395 70 -365 80
rect -215 70 -185 80
rect -20 100 50 110
rect -20 80 25 100
rect 45 80 50 100
rect -20 70 50 80
rect -890 40 -860 55
rect -710 40 -680 55
rect -530 40 -500 55
rect -350 40 -320 55
rect -170 40 -140 55
rect -890 20 -885 40
rect -865 20 -705 40
rect -685 20 -525 40
rect -505 20 -345 40
rect -325 20 -165 40
rect -145 20 -140 40
rect -890 10 -860 20
rect -710 10 -680 20
rect -530 10 -500 20
rect -350 10 -320 20
rect -170 10 -140 20
rect -20 40 10 70
rect -20 20 -15 40
rect 5 20 10 40
rect -20 10 10 20
rect 70 40 100 50
rect 70 20 75 40
rect 95 20 100 40
rect 70 -10 100 20
rect 270 40 300 50
rect 270 20 275 40
rect 295 20 300 40
rect 270 -10 300 20
rect 470 40 500 50
rect 470 20 475 40
rect 495 20 500 40
rect 470 -10 500 20
rect 670 40 700 50
rect 670 20 675 40
rect 695 20 700 40
rect 670 -10 700 20
rect 870 40 900 50
rect 870 20 875 40
rect 895 20 900 40
rect 870 -10 900 20
rect 1070 40 1100 50
rect 1070 20 1075 40
rect 1095 20 1100 40
rect 1070 -10 1100 20
rect 1270 40 1300 50
rect 1270 20 1275 40
rect 1295 20 1300 40
rect 1270 -10 1300 20
rect 1470 40 1500 50
rect 1470 20 1475 40
rect 1495 20 1500 40
rect 1470 -10 1500 20
rect 1670 40 1700 50
rect 1670 20 1675 40
rect 1695 20 1700 40
rect 1670 -10 1700 20
rect 1870 40 1900 50
rect 1870 20 1875 40
rect 1895 20 1900 40
rect 1870 -10 1900 20
rect 2070 40 2100 50
rect 2070 20 2075 40
rect 2095 20 2100 40
rect 2070 -10 2100 20
rect 2270 40 2300 50
rect 2270 20 2275 40
rect 2295 20 2300 40
rect 2270 -10 2300 20
rect 2470 40 2500 50
rect 2470 20 2475 40
rect 2495 20 2500 40
rect 2470 -10 2500 20
rect 2670 40 2700 50
rect 2670 20 2675 40
rect 2695 20 2700 40
rect 2670 -10 2700 20
rect 2790 40 2820 50
rect 2790 20 2795 40
rect 2815 20 2820 40
rect 2790 -10 2820 20
rect 70 -30 2820 -10
<< via1 >>
rect 65 150 95 155
rect 65 130 70 150
rect 70 130 90 150
rect 90 130 95 150
rect 65 125 95 130
rect 2610 125 2640 155
<< metal2 >>
rect 60 155 100 160
rect 60 125 65 155
rect 95 150 100 155
rect 2605 155 2645 160
rect 2605 150 2610 155
rect 95 130 2610 150
rect 95 125 100 130
rect 60 120 100 125
rect 2605 125 2610 130
rect 2640 125 2645 155
rect 2605 120 2645 125
use csi  csi_0
timestamp 1765329033
transform 1 0 175 0 1 0
box -125 -85 85 455
use csi  csi_1
timestamp 1765329033
transform 1 0 375 0 1 0
box -125 -85 85 455
use csi  csi_2
timestamp 1765329033
transform 1 0 575 0 1 0
box -125 -85 85 455
use csi  csi_3
timestamp 1765329033
transform 1 0 775 0 1 0
box -125 -85 85 455
use csi  csi_4
timestamp 1765329033
transform 1 0 975 0 1 0
box -125 -85 85 455
use csi  csi_5
timestamp 1765329033
transform 1 0 1175 0 1 0
box -125 -85 85 455
use csi  csi_6
timestamp 1765329033
transform 1 0 1375 0 1 0
box -125 -85 85 455
use csi  csi_7
timestamp 1765329033
transform 1 0 1575 0 1 0
box -125 -85 85 455
use csi  csi_8
timestamp 1765329033
transform 1 0 1775 0 1 0
box -125 -85 85 455
use csi  csi_9
timestamp 1765329033
transform 1 0 1975 0 1 0
box -125 -85 85 455
use csi  csi_10
timestamp 1765329033
transform 1 0 2175 0 1 0
box -125 -85 85 455
use csi  csi_11
timestamp 1765329033
transform 1 0 2375 0 1 0
box -125 -85 85 455
use csi  csi_12
timestamp 1765329033
transform 1 0 2575 0 1 0
box -125 -85 85 455
use inv  inv_0
timestamp 1765328216
transform 1 0 2690 0 1 0
box -40 -280 85 600
use inv  inv_2
timestamp 1765328216
transform 1 0 2810 0 1 0
box -40 -280 85 600
<< end >>
