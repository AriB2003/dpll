magic
tech sky130A
timestamp 1765340971
<< nwell >>
rect 290 1635 2565 1645
rect 1620 1610 2565 1635
rect 760 1585 1060 1605
rect 1600 1590 2565 1610
rect 290 1565 295 1570
rect 290 1560 300 1565
rect 290 1540 320 1560
rect 300 1415 320 1540
rect 960 1530 970 1550
rect 1620 1500 2565 1590
rect 310 1375 330 1390
rect 1750 1365 1770 1500
rect 2165 1365 2185 1500
rect 1635 1345 1665 1365
rect 2050 1345 2080 1365
rect 2165 1345 2195 1365
<< psubdiff >>
rect 2100 1145 2150 1150
rect 2100 1125 2115 1145
rect 2135 1125 2150 1145
rect 2100 1120 2150 1125
<< nsubdiff >>
rect 2100 1565 2150 1570
rect 2100 1545 2115 1565
rect 2135 1545 2150 1565
rect 2100 1540 2150 1545
<< psubdiffcont >>
rect 2115 1125 2135 1145
<< nsubdiffcont >>
rect 2115 1545 2135 1565
<< poly >>
rect 230 1530 260 1540
rect 230 1510 235 1530
rect 255 1510 260 1530
rect 230 1500 260 1510
rect 230 1495 245 1500
rect 2050 1355 2080 1365
rect 2050 1335 2055 1355
rect 2075 1335 2080 1355
rect 2050 1325 2080 1335
rect 2165 1355 2195 1365
rect 2165 1335 2170 1355
rect 2190 1335 2195 1355
rect 2165 1325 2195 1335
rect 230 1190 245 1195
rect 230 1180 260 1190
rect 230 1160 235 1180
rect 255 1160 260 1180
rect 230 1150 260 1160
<< polycont >>
rect 235 1510 255 1530
rect 2055 1335 2075 1355
rect 2170 1335 2190 1355
rect 235 1160 255 1180
<< locali >>
rect 230 1590 285 1610
rect 265 1575 285 1590
rect 1890 1580 2075 1600
rect 2305 1580 2490 1600
rect 265 1570 290 1575
rect 265 1565 295 1570
rect 265 1560 300 1565
rect 270 1555 320 1560
rect 275 1550 320 1555
rect 280 1540 320 1550
rect 230 1530 260 1540
rect 230 1510 235 1530
rect 255 1510 260 1530
rect 230 1500 260 1510
rect 300 1430 320 1540
rect 2055 1515 2075 1580
rect 2105 1565 2145 1570
rect 2105 1545 2115 1565
rect 2135 1545 2145 1565
rect 2105 1540 2145 1545
rect 2115 1515 2135 1540
rect 2470 1515 2490 1580
rect 300 1420 330 1430
rect 300 1400 305 1420
rect 325 1400 330 1420
rect 300 1390 330 1400
rect 1635 1355 1665 1365
rect 280 1335 350 1355
rect 930 1335 1010 1355
rect 1635 1335 1640 1355
rect 1660 1335 1665 1355
rect 1635 1325 1665 1335
rect 1750 1355 1780 1365
rect 1750 1335 1755 1355
rect 1775 1335 1780 1355
rect 1750 1325 1780 1335
rect 2050 1355 2080 1365
rect 2050 1335 2055 1355
rect 2075 1335 2080 1355
rect 2050 1325 2080 1335
rect 2165 1355 2195 1365
rect 2165 1335 2170 1355
rect 2190 1335 2195 1355
rect 2430 1335 2460 1355
rect 2165 1325 2195 1335
rect 190 1210 200 1260
rect 190 1110 210 1210
rect 230 1180 260 1190
rect 230 1160 235 1180
rect 255 1160 260 1180
rect 230 1150 260 1160
rect 1640 1115 1660 1175
rect 2115 1150 2135 1175
rect 2105 1145 2145 1150
rect 2105 1125 2115 1145
rect 2135 1125 2145 1145
rect 2105 1120 2145 1125
rect 190 1100 225 1110
rect 190 1080 200 1100
rect 220 1080 225 1100
rect 190 1070 225 1080
rect 1640 1105 1670 1115
rect 1640 1085 1645 1105
rect 1665 1085 1670 1105
rect 2200 1110 2230 1120
rect 2200 1100 2205 1110
rect 1640 1075 1670 1085
rect 2015 1090 2205 1100
rect 2225 1090 2230 1110
rect 2015 1080 2230 1090
rect 2265 1065 2285 1070
rect 1870 1060 1890 1065
rect 2265 1060 2305 1065
rect 2470 1060 2490 1175
rect 1870 1040 2490 1060
<< viali >>
rect 1865 1590 1885 1610
rect 235 1510 255 1530
rect 200 1445 220 1465
rect 305 1400 325 1420
rect 1640 1335 1660 1355
rect 1755 1335 1775 1355
rect 2055 1335 2075 1355
rect 2170 1335 2190 1355
rect 235 1160 255 1180
rect 200 1080 220 1100
rect 1645 1085 1665 1105
rect 2205 1090 2225 1110
<< metal1 >>
rect 270 1635 2185 1655
rect 270 1550 290 1635
rect 1860 1610 1890 1620
rect 760 1585 1060 1605
rect 1600 1590 1865 1610
rect 1885 1590 1890 1610
rect 1860 1580 1890 1590
rect 230 1530 310 1550
rect 960 1530 970 1550
rect 1620 1530 1770 1550
rect 230 1510 235 1530
rect 255 1510 260 1530
rect 230 1500 260 1510
rect 195 1470 225 1475
rect 195 1435 225 1440
rect 300 1420 330 1430
rect 300 1400 305 1420
rect 325 1400 330 1420
rect 300 1390 330 1400
rect 310 1355 330 1390
rect 1750 1365 1770 1530
rect 2165 1365 2185 1635
rect 1635 1355 1665 1365
rect 310 1335 350 1355
rect 930 1335 1010 1355
rect 1635 1335 1640 1355
rect 1660 1335 1665 1355
rect 1635 1325 1665 1335
rect 1750 1355 1780 1365
rect 1750 1335 1755 1355
rect 1775 1335 1780 1355
rect 1750 1325 1780 1335
rect 2050 1355 2080 1365
rect 2050 1335 2055 1355
rect 2075 1335 2080 1355
rect 2050 1325 2080 1335
rect 2165 1355 2195 1365
rect 2165 1335 2170 1355
rect 2190 1335 2195 1355
rect 2165 1325 2195 1335
rect 230 1180 260 1190
rect 230 1160 235 1180
rect 255 1160 260 1180
rect 230 1140 310 1160
rect 960 1140 970 1160
rect 195 1100 225 1110
rect 195 1080 200 1100
rect 220 1080 225 1100
rect 940 1080 970 1100
rect 195 1070 225 1080
rect 1020 1055 1040 1160
rect 1645 1155 1665 1325
rect 1645 1135 1710 1155
rect 1640 1105 1670 1115
rect 1420 1085 1645 1105
rect 1665 1085 1670 1105
rect 1640 1075 1670 1085
rect 1690 1055 1710 1135
rect 2050 1055 2070 1325
rect 2200 1110 2230 1120
rect 2200 1090 2205 1110
rect 2225 1100 2230 1110
rect 2225 1090 2545 1100
rect 2200 1080 2545 1090
rect 1020 1035 2070 1055
<< via1 >>
rect 195 1465 225 1470
rect 195 1445 200 1465
rect 200 1445 220 1465
rect 220 1445 225 1465
rect 195 1440 225 1445
<< metal2 >>
rect 200 1475 220 1590
rect 190 1470 230 1475
rect 190 1440 195 1470
rect 225 1440 230 1470
rect 190 1435 230 1440
use inv  inv_0
timestamp 1765330272
transform 1 0 215 0 1 1205
box -40 -10 85 295
use inv  inv_1
timestamp 1765330272
transform 1 0 2480 0 1 1205
box -40 -10 85 295
use negdff  negdff_0
timestamp 1765332816
transform 1 0 1205 0 1 1110
box -255 -75 415 545
use posdff  posdff_0
timestamp 1765332816
transform 1 0 875 0 1 1110
box -585 -75 85 545
use xor  xor_0
timestamp 1765331190
transform 1 0 1950 0 1 1205
box -340 -155 85 440
use xor  xor_1
timestamp 1765331190
transform 1 0 2365 0 1 1205
box -340 -155 85 440
<< end >>
