magic
tech sky130A
timestamp 1765325780
<< error_s >>
rect -2942 640 -2820 645
rect -2815 615 -2725 640
rect -2815 545 -2693 615
<< nwell >>
rect 3735 545 3880 640
rect -4410 470 -2755 490
rect -4410 305 -4390 470
rect -2785 425 -2755 470
rect -480 220 -430 240
rect -25 220 10 240
rect -480 200 -460 220
<< locali >>
rect -2785 455 -2755 465
rect -2785 435 -2780 455
rect -2760 435 -2755 455
rect -2785 425 -2755 435
rect -480 220 -430 240
rect -25 220 10 240
rect -480 200 -460 220
rect -430 140 -390 145
rect -430 120 -420 140
rect -400 120 -390 140
rect -430 115 -390 120
<< viali >>
rect -2780 435 -2760 455
rect -420 120 -400 140
<< metal1 >>
rect -4410 470 -2755 490
rect -4410 305 -4390 470
rect -2785 455 -2755 470
rect -2785 435 -2780 455
rect -2760 435 -2755 455
rect -2785 425 -2755 435
rect -30 170 965 190
rect -430 140 -390 145
rect -430 120 -420 140
rect -400 120 -390 140
rect -75 120 50 140
rect -430 115 -390 120
rect -430 -65 -410 115
rect -460 -85 -410 -65
use div8  div8_0
timestamp 1765325266
transform 1 0 -5895 0 1 -260
box 700 40 3075 905
use hpd  hpd_0
timestamp 1765325701
transform 1 0 -3005 0 1 -1165
box 175 945 2565 1810
use ipump  ipump_0
timestamp 1765147879
transform 1 0 -90 0 1 40
box -360 -80 85 400
use vco  vco_0
timestamp 1765262567
transform 1 0 985 0 1 40
box -1000 -220 2895 600
<< end >>
