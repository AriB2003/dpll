magic
tech sky130A
timestamp 1765333169
<< nwell >>
rect 100 520 120 575
rect 100 500 655 520
rect 50 455 80 470
rect 85 440 180 460
rect 160 420 180 440
rect 50 390 95 410
<< locali >>
rect 50 460 80 470
rect 50 440 55 460
rect 75 440 80 460
rect 50 430 80 440
rect 55 370 75 430
rect 160 420 180 440
rect 125 380 130 420
rect 680 390 720 410
rect 50 360 80 370
rect 50 340 55 360
rect 75 340 80 360
rect 50 330 80 340
rect 110 355 130 380
rect 220 355 260 360
rect 110 335 230 355
rect 250 335 260 355
rect 220 330 260 335
<< viali >>
rect 665 500 685 520
rect 55 440 75 460
rect 55 340 75 360
rect 230 335 250 355
<< metal1 >>
rect 60 470 80 605
rect 660 525 690 530
rect 660 490 690 495
rect 50 460 80 470
rect 50 440 55 460
rect 75 440 80 460
rect 50 430 80 440
rect 50 390 95 410
rect 50 360 80 370
rect 50 340 55 360
rect 75 340 80 360
rect 50 330 80 340
rect 220 330 225 360
rect 255 330 260 360
rect 60 215 80 330
<< via1 >>
rect 95 580 125 610
rect 660 520 690 525
rect 660 500 665 520
rect 665 500 685 520
rect 685 500 690 520
rect 660 495 690 500
rect 225 355 255 360
rect 225 335 230 355
rect 230 335 250 355
rect 250 335 255 355
rect 225 330 255 335
rect 610 335 640 365
<< metal2 >>
rect 90 610 130 615
rect 90 580 95 610
rect 125 580 130 610
rect 90 575 130 580
rect 100 520 120 575
rect 655 525 695 530
rect 655 520 660 525
rect 100 500 660 520
rect 655 495 660 500
rect 690 495 695 525
rect 655 490 695 495
rect 605 365 645 370
rect 220 360 260 365
rect 605 360 610 365
rect 220 330 225 360
rect 255 335 610 360
rect 640 335 645 365
rect 255 330 260 335
rect 605 330 645 335
rect 220 325 260 330
use inv  inv_0
timestamp 1765330272
transform 1 0 740 0 1 260
box -40 -10 85 295
use posdff  posdff_0
timestamp 1765332816
transform 1 0 625 0 1 165
box -585 -75 85 545
<< end >>
