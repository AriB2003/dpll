magic
tech sky130A
timestamp 1765346501
<< error_p >>
rect -125 140 85 295
rect -10 55 15 105
rect -105 5 -70 55
rect -20 5 15 55
rect 30 55 55 105
rect 30 5 65 55
<< nwell >>
rect -125 140 85 295
<< nmos >>
rect -70 5 -20 55
rect 15 5 30 105
<< pmos >>
rect -70 225 -20 275
rect 15 175 30 275
<< ndiff >>
rect -10 55 15 105
rect -105 40 -70 55
rect -105 20 -100 40
rect -80 20 -70 40
rect -105 5 -70 20
rect -20 5 15 55
rect 30 55 55 105
rect 30 40 65 55
rect 30 20 40 40
rect 60 20 65 40
rect 30 5 65 20
<< pdiff >>
rect -105 260 -70 275
rect -105 240 -100 260
rect -80 240 -70 260
rect -105 225 -70 240
rect -20 225 15 275
rect -10 175 15 225
rect 30 260 65 275
rect 30 240 40 260
rect 60 240 65 260
rect 30 225 65 240
rect 30 175 55 225
<< ndiffc >>
rect -100 20 -80 40
rect 40 20 60 40
<< pdiffc >>
rect -100 240 -80 260
rect 40 240 60 260
<< poly >>
rect -70 275 -20 290
rect 15 275 30 290
rect -70 210 -20 225
rect -65 200 -35 210
rect -65 180 -60 200
rect -40 180 -35 200
rect -65 170 -35 180
rect 15 160 30 175
rect -15 150 30 160
rect -15 130 -10 150
rect 10 130 30 150
rect -15 120 30 130
rect -65 100 -35 110
rect 15 105 30 120
rect -65 80 -60 100
rect -40 80 -35 100
rect -65 70 -35 80
rect -70 55 -20 70
rect -70 -10 -20 5
rect 15 -10 30 5
<< polycont >>
rect -60 180 -40 200
rect -10 130 10 150
rect -60 80 -40 100
<< locali >>
rect -105 260 -75 275
rect -105 240 -100 260
rect -80 240 -75 260
rect -105 225 -75 240
rect 35 260 65 270
rect 35 240 40 260
rect 60 240 65 260
rect 35 225 65 240
rect -65 200 -35 210
rect -105 180 -60 200
rect -40 180 65 200
rect -65 170 -35 180
rect -15 150 15 160
rect -105 130 -10 150
rect 10 130 15 150
rect -15 120 15 130
rect 35 150 65 160
rect 35 130 40 150
rect 60 130 65 150
rect 35 120 65 130
rect -65 100 -35 110
rect -105 80 -60 100
rect -40 80 65 100
rect -65 70 -35 80
rect -105 40 -75 55
rect -105 20 -100 40
rect -80 20 -75 40
rect -105 5 -75 20
rect 35 40 65 55
rect 35 20 40 40
rect 60 20 65 40
rect 35 10 65 20
<< viali >>
rect 40 240 60 260
rect 40 130 60 150
rect 40 20 60 40
<< metal1 >>
rect 35 260 65 270
rect 35 240 40 260
rect 60 240 65 260
rect 35 150 65 240
rect 35 130 40 150
rect 60 130 65 150
rect 35 40 65 130
rect 35 20 40 40
rect 60 20 65 40
rect 35 10 65 20
<< end >>
