magic
tech sky130A
timestamp 1765329072
<< nwell >>
rect 270 1655 290 1660
rect 840 1655 1095 1810
rect 1960 1730 2115 1810
rect 2310 1710 2565 1810
rect 270 1635 2185 1655
rect 270 1610 290 1635
rect 1860 1610 1890 1620
rect 230 1590 290 1610
rect 265 1570 290 1590
rect 760 1585 1060 1605
rect 1600 1600 1890 1610
rect 1600 1590 2075 1600
rect 1860 1580 2075 1590
rect 265 1565 295 1570
rect 265 1560 300 1565
rect 270 1550 320 1560
rect 280 1540 320 1550
rect 300 1415 320 1540
rect 960 1530 970 1550
rect 1620 1530 1770 1550
rect 1750 1365 1770 1530
rect 2055 1515 2075 1580
rect 2165 1365 2185 1635
rect 2305 1580 2490 1600
rect 2470 1515 2490 1580
rect 1635 1345 1665 1365
rect 2050 1345 2080 1365
rect 2165 1345 2195 1365
<< poly >>
rect 230 1530 260 1540
rect 230 1510 235 1530
rect 255 1510 260 1530
rect 230 1500 260 1510
rect 230 1495 245 1500
rect 2050 1355 2080 1365
rect 2050 1335 2055 1355
rect 2075 1335 2080 1355
rect 2050 1325 2080 1335
rect 2165 1355 2195 1365
rect 2165 1335 2170 1355
rect 2190 1335 2195 1355
rect 2165 1325 2195 1335
rect 230 1190 245 1195
rect 230 1180 260 1190
rect 230 1160 235 1180
rect 255 1160 260 1180
rect 230 1150 260 1160
<< polycont >>
rect 235 1510 255 1530
rect 2055 1335 2075 1355
rect 2170 1335 2190 1355
rect 235 1160 255 1180
<< locali >>
rect 230 1590 285 1610
rect 265 1575 285 1590
rect 1890 1580 2075 1600
rect 2305 1580 2490 1600
rect 265 1570 290 1575
rect 265 1565 295 1570
rect 265 1560 300 1565
rect 270 1555 320 1560
rect 275 1550 320 1555
rect 280 1540 320 1550
rect 230 1530 260 1540
rect 230 1510 235 1530
rect 255 1510 260 1530
rect 230 1500 260 1510
rect 300 1415 320 1540
rect 2055 1515 2075 1580
rect 2470 1515 2490 1580
rect 300 1405 330 1415
rect 300 1385 305 1405
rect 325 1385 330 1405
rect 300 1375 330 1385
rect 1635 1355 1665 1365
rect 280 1335 350 1355
rect 930 1335 1010 1355
rect 1635 1335 1640 1355
rect 1660 1335 1665 1355
rect 1635 1325 1665 1335
rect 1750 1355 1780 1365
rect 1750 1335 1755 1355
rect 1775 1335 1780 1355
rect 1750 1325 1780 1335
rect 2050 1355 2080 1365
rect 2050 1335 2055 1355
rect 2075 1335 2080 1355
rect 2050 1325 2080 1335
rect 2165 1355 2195 1365
rect 2165 1335 2170 1355
rect 2190 1335 2195 1355
rect 2430 1335 2460 1355
rect 2165 1325 2195 1335
rect 230 1180 260 1190
rect 230 1160 235 1180
rect 255 1160 260 1180
rect 230 1150 260 1160
rect 1640 1115 1660 1175
rect 1640 1105 1670 1115
rect 1640 1085 1645 1105
rect 1665 1085 1670 1105
rect 2095 1110 2125 1120
rect 2095 1100 2100 1110
rect 1640 1075 1670 1085
rect 2015 1090 2100 1100
rect 2120 1090 2125 1110
rect 2015 1080 2125 1090
rect 2265 1065 2285 1070
rect 1870 1060 1890 1065
rect 2265 1060 2305 1065
rect 2470 1060 2490 1175
rect 1870 1040 2490 1060
<< viali >>
rect 1865 1590 1885 1610
rect 235 1510 255 1530
rect 305 1385 325 1405
rect 1640 1335 1660 1355
rect 1755 1335 1775 1355
rect 2055 1335 2075 1355
rect 2170 1335 2190 1355
rect 235 1160 255 1180
rect 1645 1085 1665 1105
rect 2100 1090 2120 1110
<< metal1 >>
rect 270 1635 2185 1655
rect 270 1550 290 1635
rect 1860 1610 1890 1620
rect 760 1585 1060 1605
rect 1600 1590 1865 1610
rect 1885 1590 1890 1610
rect 1860 1580 1890 1590
rect 230 1530 310 1550
rect 960 1530 970 1550
rect 1620 1530 1770 1550
rect 230 1510 235 1530
rect 255 1510 260 1530
rect 230 1500 260 1510
rect 300 1405 330 1415
rect 300 1385 305 1405
rect 325 1385 330 1405
rect 300 1375 330 1385
rect 310 1355 330 1375
rect 1750 1365 1770 1530
rect 2165 1365 2185 1635
rect 1635 1355 1665 1365
rect 310 1335 350 1355
rect 930 1335 1010 1355
rect 1635 1335 1640 1355
rect 1660 1335 1665 1355
rect 1635 1325 1665 1335
rect 1750 1355 1780 1365
rect 1750 1335 1755 1355
rect 1775 1335 1780 1355
rect 1750 1325 1780 1335
rect 2050 1355 2080 1365
rect 2050 1335 2055 1355
rect 2075 1335 2080 1355
rect 2050 1325 2080 1335
rect 2165 1355 2195 1365
rect 2165 1335 2170 1355
rect 2190 1335 2195 1355
rect 2165 1325 2195 1335
rect 230 1180 260 1190
rect 230 1160 235 1180
rect 255 1160 260 1180
rect 230 1140 310 1160
rect 960 1140 970 1160
rect 940 1080 970 1100
rect 1020 1055 1040 1160
rect 1645 1155 1665 1325
rect 1645 1135 1710 1155
rect 1640 1105 1670 1115
rect 1420 1085 1645 1105
rect 1665 1085 1670 1105
rect 1640 1075 1670 1085
rect 1690 1055 1710 1135
rect 2050 1055 2070 1325
rect 2095 1110 2125 1120
rect 2095 1090 2100 1110
rect 2120 1100 2125 1110
rect 2120 1090 2545 1100
rect 2095 1080 2545 1090
rect 1020 1035 2070 1055
use inv  inv_0
timestamp 1765328216
transform 1 0 215 0 1 1205
box -40 -280 85 600
use inv  inv_1
timestamp 1765328216
transform 1 0 2480 0 1 1205
box -40 -280 85 600
use negdff  negdff_0
timestamp 1765307306
transform 1 0 1205 0 1 1110
box -295 -165 415 700
use posdff  posdff_0
timestamp 1765307294
transform 1 0 875 0 1 1110
box -625 -165 85 700
use xor  xor_0
timestamp 1765328216
transform 1 0 1950 0 1 1205
box -340 -280 85 605
use xor  xor_1
timestamp 1765328216
transform 1 0 2365 0 1 1205
box -340 -280 85 605
<< end >>
