magic
tech sky130A
timestamp 1765307306
<< nwell >>
rect -115 480 95 500
rect 85 420 95 440
<< locali >>
rect 55 225 135 245
<< metal1 >>
rect -115 480 95 500
rect 85 420 95 440
rect 55 225 135 245
rect 85 30 95 50
rect 65 -30 185 -10
use csrl  csrl_0
timestamp 1765307270
transform 1 0 330 0 1 30
box -295 -165 85 640
use ncsrl  ncsrl_0
timestamp 1765307252
transform 1 0 0 0 1 95
box -295 -260 85 605
<< end >>
