magic
tech sky130A
timestamp 1765406647
<< locali >>
rect -4430 485 -4390 490
rect -4430 465 -4420 485
rect -4400 465 -4390 485
rect -4430 460 -4390 465
rect -5130 425 -5110 445
rect -4410 310 -4390 460
rect -2785 455 -2755 465
rect -2785 435 -2780 455
rect -2760 435 -2755 455
rect -2785 425 -2755 435
rect -535 330 -410 350
rect -535 315 -515 330
rect -430 315 -410 330
rect -25 220 10 240
rect -2800 170 -2780 190
rect 3835 170 3855 190
rect -50 60 -30 80
rect 100 60 120 80
rect -535 30 -515 45
rect -430 30 -410 45
rect -535 10 -410 30
rect -5040 -80 -5020 -60
<< viali >>
rect -4420 465 -4400 485
rect -2780 435 -2760 455
<< metal1 >>
rect -4430 485 -2755 490
rect -4430 465 -4420 485
rect -4400 470 -2755 485
rect -4400 465 -4390 470
rect -4430 460 -4390 465
rect -2785 455 -2755 470
rect -2925 450 -2895 455
rect -2785 435 -2780 455
rect -2760 435 -2755 455
rect -2785 425 -2755 435
rect -2925 415 -2895 420
rect -430 330 125 350
rect 95 315 125 330
rect -4410 305 -4390 310
rect -460 195 -430 225
rect -30 170 965 190
rect -430 -65 -410 135
rect -75 120 50 140
rect -385 10 1055 30
rect -2955 -85 -2605 -65
rect -460 -85 -410 -65
<< via1 >>
rect -3165 415 -3135 445
rect -2925 420 -2895 450
rect -2695 420 -2665 450
rect -4995 165 -4965 195
rect 3830 165 3860 195
<< metal2 >>
rect -2930 450 -2890 455
rect -3170 445 -3130 450
rect -2930 445 -2925 450
rect -3170 415 -3165 445
rect -3135 425 -2925 445
rect -3135 415 -3130 425
rect -2930 420 -2925 425
rect -2895 445 -2890 450
rect -2700 450 -2660 455
rect -2700 445 -2695 450
rect -2895 425 -2695 445
rect -2895 420 -2890 425
rect -2930 415 -2890 420
rect -2700 420 -2695 425
rect -2665 420 -2660 450
rect -2700 415 -2660 420
rect -3170 410 -3130 415
rect -4995 230 3865 250
rect -4995 200 -4970 230
rect -5000 195 -4960 200
rect -5000 165 -4995 195
rect -4965 165 -4960 195
rect -5000 160 -4960 165
rect 3825 195 3865 230
rect 3825 165 3830 195
rect 3860 165 3865 195
rect 3825 160 3865 165
use div8  div8_0
timestamp 1765346567
transform 1 0 -5895 0 1 -260
box 740 130 3075 750
use hpd  hpd_0
timestamp 1765346567
transform 1 0 -3005 0 1 -1165
box 175 1035 2565 1655
use ipump  ipump_0
timestamp 1765330714
transform 1 0 -90 0 1 40
box -360 -25 85 300
use vco  vco_0
timestamp 1765346501
transform 1 0 985 0 1 40
box -1000 -55 2895 355
<< labels >>
rlabel via1 3845 180 3845 180 3 clk
port 4 e
rlabel locali -5120 435 -5120 435 7 VP
port 1 w
rlabel locali -5030 -70 -5030 -70 7 VN
port 2 w
rlabel locali -2790 180 -2790 180 7 nrz
port 3 w
rlabel locali 110 70 110 70 7 res
port 5 w
rlabel locali -40 70 -40 70 7 filt
port 6 w
<< end >>
