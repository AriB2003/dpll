* SPICE3 file created from dpll.ext - technology: sky130A

X0 m1_n8820_610# div8_0/div_0/li_100_660# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.175 ps=1.7 w=0.5 l=0.15
X1 m1_n8820_610# div8_0/div_0/li_100_660# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.175 ps=1.7 w=0.5 l=0.15
X2 div8_0/div_0/posdff_0/li_n550_450# div8_0/div_0/posdff_0/m1_n490_60# div8_0/div_0/posdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.1 ps=0.9 w=0.5 l=0.5
X3 div8_0/div_0/posdff_0/csrl_0/a_n470_n150# m1_n9990_330# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1475 ps=1.275 w=0.5 l=0.5
X4 div8_0/div_0/posdff_0/csrl_0/a_n300_580# div8_0/div_0/li_220_670# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.24625 ps=2.5 w=0.5 l=0.5
X5 div8_0/div_0/posdff_0/csrl_0/a_n470_140# m1_n9990_330# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1475 ps=1.275 w=0.5 l=0.5
X6 m1_n860_660# div8_0/div_0/posdff_0/m1_n490_60# div8_0/div_0/posdff_0/li_n550_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.24625 pd=2.5 as=0.1 ps=0.9 w=0.5 l=0.5
X7 VSUBS div8_0/div_0/li_100_660# div8_0/div_0/posdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.19665 pd=1.7 as=0.175 ps=1.7 w=0.5 l=0.5
X8 div8_0/div_0/posdff_0/li_n550_450# m1_n9990_330# div8_0/div_0/posdff_0/csrl_0/a_n300_580# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X9 div8_0/div_0/posdff_0/csrl_0/a_n300_870# div8_0/div_0/li_100_660# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.24625 ps=2.5 w=0.5 l=0.5
X10 div8_0/div_0/posdff_0/m1_n490_60# div8_0/div_0/posdff_0/li_n550_450# div8_0/div_0/posdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.1 ps=0.9 w=0.5 l=0.5
X11 m1_n860_660# div8_0/div_0/posdff_0/li_n550_450# div8_0/div_0/posdff_0/m1_n490_60# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.24625 pd=2.5 as=0.1 ps=0.9 w=0.5 l=0.5
X12 VSUBS div8_0/div_0/li_220_670# div8_0/div_0/posdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0.19665 pd=1.7 as=0.175 ps=1.7 w=0.5 l=0.5
X13 div8_0/div_0/posdff_0/m1_n490_60# m1_n9990_330# div8_0/div_0/posdff_0/csrl_0/a_n300_870# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X14 div8_0/div_0/li_220_670# div8_0/div_0/li_100_660# div8_0/div_0/posdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.1 ps=0.9 w=0.5 l=0.5
X15 div8_0/div_0/posdff_0/ncsrl_0/a_n470_740# m1_n9990_330# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1475 ps=1.275 w=0.5 l=0.5
X16 div8_0/div_0/li_100_660# m1_n9990_330# div8_0/div_0/posdff_0/ncsrl_0/a_n300_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X17 div8_0/div_0/posdff_0/ncsrl_0/a_n300_n280# div8_0/div_0/posdff_0/m1_n490_60# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.24625 ps=2.5 w=0.5 l=0.5
X18 VSUBS div8_0/div_0/li_220_670# div8_0/div_0/li_100_660# VSUBS sky130_fd_pr__nfet_01v8 ad=0.24625 pd=2.5 as=0.1 ps=0.9 w=0.5 l=0.5
X19 div8_0/div_0/posdff_0/ncsrl_0/a_n300_10# div8_0/div_0/posdff_0/li_n550_450# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.24625 ps=2.5 w=0.5 l=0.5
X20 m1_n860_660# div8_0/div_0/posdff_0/li_n550_450# div8_0/div_0/posdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.19665 pd=1.7 as=0.175 ps=1.7 w=0.5 l=0.5
X21 VSUBS div8_0/div_0/li_100_660# div8_0/div_0/li_220_670# VSUBS sky130_fd_pr__nfet_01v8 ad=0.24625 pd=2.5 as=0.1 ps=0.9 w=0.5 l=0.5
X22 div8_0/div_0/li_100_660# div8_0/div_0/li_220_670# div8_0/div_0/posdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.1 ps=0.9 w=0.5 l=0.5
X23 div8_0/div_0/posdff_0/ncsrl_0/a_n470_450# m1_n9990_330# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1475 ps=1.275 w=0.5 l=0.5
X24 m1_n860_660# div8_0/div_0/posdff_0/m1_n490_60# div8_0/div_0/posdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.19665 pd=1.7 as=0.175 ps=1.7 w=0.5 l=0.5
X25 div8_0/div_0/li_220_670# m1_n9990_330# div8_0/div_0/posdff_0/ncsrl_0/a_n300_n280# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X26 div8_0/m1_4560_860# div8_0/div_1/li_100_660# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=13.46 ps=128.905 w=0.5 l=0.15
X27 div8_0/m1_4560_860# div8_0/div_1/li_100_660# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=14.46 ps=137.905 w=0.5 l=0.15
X28 div8_0/div_1/posdff_0/li_n550_450# div8_0/div_1/posdff_0/m1_n490_60# div8_0/div_1/posdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.375 ps=3.5 w=0.5 l=0.5
X29 div8_0/div_1/posdff_0/csrl_0/a_n470_n150# m1_n8820_610# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.375 pd=3.5 as=0 ps=0 w=0.5 l=0.5
X30 div8_0/div_1/posdff_0/csrl_0/a_n300_580# div8_0/div_1/li_220_670# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X31 div8_0/div_1/posdff_0/csrl_0/a_n470_140# m1_n8820_610# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X32 m1_n860_660# div8_0/div_1/posdff_0/m1_n490_60# div8_0/div_1/posdff_0/li_n550_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X33 VSUBS div8_0/div_1/li_100_660# div8_0/div_1/posdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X34 div8_0/div_1/posdff_0/li_n550_450# m1_n8820_610# div8_0/div_1/posdff_0/csrl_0/a_n300_580# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X35 div8_0/div_1/posdff_0/csrl_0/a_n300_870# div8_0/div_1/li_100_660# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X36 div8_0/div_1/posdff_0/m1_n490_60# div8_0/div_1/posdff_0/li_n550_450# div8_0/div_1/posdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.5
X37 m1_n860_660# div8_0/div_1/posdff_0/li_n550_450# div8_0/div_1/posdff_0/m1_n490_60# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X38 VSUBS div8_0/div_1/li_220_670# div8_0/div_1/posdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X39 div8_0/div_1/posdff_0/m1_n490_60# m1_n8820_610# div8_0/div_1/posdff_0/csrl_0/a_n300_870# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X40 div8_0/div_1/li_220_670# div8_0/div_1/li_100_660# div8_0/div_1/posdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.375 ps=3.5 w=0.5 l=0.5
X41 div8_0/div_1/posdff_0/ncsrl_0/a_n470_740# m1_n8820_610# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X42 div8_0/div_1/li_100_660# m1_n8820_610# div8_0/div_1/posdff_0/ncsrl_0/a_n300_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.5
X43 div8_0/div_1/posdff_0/ncsrl_0/a_n300_n280# div8_0/div_1/posdff_0/m1_n490_60# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X44 VSUBS div8_0/div_1/li_220_670# div8_0/div_1/li_100_660# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X45 div8_0/div_1/posdff_0/ncsrl_0/a_n300_10# div8_0/div_1/posdff_0/li_n550_450# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X46 m1_n860_660# div8_0/div_1/posdff_0/li_n550_450# div8_0/div_1/posdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.375 ps=3.5 w=0.5 l=0.5
X47 VSUBS div8_0/div_1/li_100_660# div8_0/div_1/li_220_670# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X48 div8_0/div_1/li_100_660# div8_0/div_1/li_220_670# div8_0/div_1/posdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.5
X49 div8_0/div_1/posdff_0/ncsrl_0/a_n470_450# m1_n8820_610# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X50 m1_n860_660# div8_0/div_1/posdff_0/m1_n490_60# div8_0/div_1/posdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X51 div8_0/div_1/li_220_670# m1_n8820_610# div8_0/div_1/posdff_0/ncsrl_0/a_n300_n280# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X52 div8_0/div_2/inv_0/a_60_10# div8_0/div_2/li_100_660# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X53 div8_0/div_2/inv_0/a_60_10# div8_0/div_2/li_100_660# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X54 div8_0/div_2/posdff_0/li_n550_450# div8_0/div_2/posdff_0/m1_n490_60# div8_0/div_2/posdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.375 ps=3.5 w=0.5 l=0.5
X55 div8_0/div_2/posdff_0/csrl_0/a_n470_n150# div8_0/m1_4560_860# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.375 pd=3.5 as=0 ps=0 w=0.5 l=0.5
X56 div8_0/div_2/posdff_0/csrl_0/a_n300_580# div8_0/div_2/li_220_670# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X57 div8_0/div_2/posdff_0/csrl_0/a_n470_140# div8_0/m1_4560_860# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X58 m1_n860_660# div8_0/div_2/posdff_0/m1_n490_60# div8_0/div_2/posdff_0/li_n550_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X59 VSUBS div8_0/div_2/li_100_660# div8_0/div_2/posdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X60 div8_0/div_2/posdff_0/li_n550_450# div8_0/m1_4560_860# div8_0/div_2/posdff_0/csrl_0/a_n300_580# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X61 div8_0/div_2/posdff_0/csrl_0/a_n300_870# div8_0/div_2/li_100_660# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X62 div8_0/div_2/posdff_0/m1_n490_60# div8_0/div_2/posdff_0/li_n550_450# div8_0/div_2/posdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.5
X63 m1_n860_660# div8_0/div_2/posdff_0/li_n550_450# div8_0/div_2/posdff_0/m1_n490_60# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X64 VSUBS div8_0/div_2/li_220_670# div8_0/div_2/posdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X65 div8_0/div_2/posdff_0/m1_n490_60# div8_0/m1_4560_860# div8_0/div_2/posdff_0/csrl_0/a_n300_870# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X66 div8_0/div_2/li_220_670# div8_0/div_2/li_100_660# div8_0/div_2/posdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.375 ps=3.5 w=0.5 l=0.5
X67 div8_0/div_2/posdff_0/ncsrl_0/a_n470_740# div8_0/m1_4560_860# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X68 div8_0/div_2/li_100_660# div8_0/m1_4560_860# div8_0/div_2/posdff_0/ncsrl_0/a_n300_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.5
X69 div8_0/div_2/posdff_0/ncsrl_0/a_n300_n280# div8_0/div_2/posdff_0/m1_n490_60# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X70 VSUBS div8_0/div_2/li_220_670# div8_0/div_2/li_100_660# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X71 div8_0/div_2/posdff_0/ncsrl_0/a_n300_10# div8_0/div_2/posdff_0/li_n550_450# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X72 m1_n860_660# div8_0/div_2/posdff_0/li_n550_450# div8_0/div_2/posdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.375 ps=3.5 w=0.5 l=0.5
X73 VSUBS div8_0/div_2/li_100_660# div8_0/div_2/li_220_670# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X74 div8_0/div_2/li_100_660# div8_0/div_2/li_220_670# div8_0/div_2/posdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.5
X75 div8_0/div_2/posdff_0/ncsrl_0/a_n470_450# div8_0/m1_4560_860# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X76 m1_n860_660# div8_0/div_2/posdff_0/m1_n490_60# div8_0/div_2/posdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X77 div8_0/div_2/li_220_670# div8_0/m1_4560_860# div8_0/div_2/posdff_0/ncsrl_0/a_n300_n280# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X78 hpd_0/negdff_0/csrl_0/a_n120_580# hpd_0/li_3500_2650# hpd_0/negdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.375 ps=3.5 w=0.5 l=0.5
X79 hpd_0/negdff_0/csrl_0/a_n470_n150# m1_n8820_610# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.375 pd=3.5 as=0 ps=0 w=0.5 l=0.5
X80 hpd_0/negdff_0/csrl_0/a_n300_580# hpd_0/negdff_0/li_110_450# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X81 hpd_0/negdff_0/csrl_0/a_n470_140# m1_n8820_610# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X82 m1_n860_660# hpd_0/li_3500_2650# hpd_0/negdff_0/csrl_0/a_n120_580# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X83 VSUBS hpd_0/negdff_0/m1_170_60# hpd_0/negdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X84 hpd_0/negdff_0/csrl_0/a_n120_580# m1_n8820_610# hpd_0/negdff_0/csrl_0/a_n300_580# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X85 hpd_0/negdff_0/csrl_0/a_n300_870# hpd_0/negdff_0/m1_170_60# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X86 hpd_0/li_3500_2650# hpd_0/negdff_0/csrl_0/a_n120_580# hpd_0/negdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.5
X87 m1_n860_660# hpd_0/negdff_0/csrl_0/a_n120_580# hpd_0/li_3500_2650# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X88 VSUBS hpd_0/negdff_0/li_110_450# hpd_0/negdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X89 hpd_0/li_3500_2650# m1_n8820_610# hpd_0/negdff_0/csrl_0/a_n300_870# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X90 hpd_0/negdff_0/m1_170_60# hpd_0/negdff_0/li_110_450# hpd_0/negdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.375 ps=3.5 w=0.5 l=0.5
X91 hpd_0/negdff_0/ncsrl_0/a_n470_740# m1_n8820_610# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X92 hpd_0/negdff_0/li_110_450# m1_n8820_610# hpd_0/negdff_0/ncsrl_0/a_n300_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.5
X93 hpd_0/negdff_0/ncsrl_0/a_n300_n280# hpd_0/a_4100_2650# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X94 VSUBS hpd_0/negdff_0/m1_170_60# hpd_0/negdff_0/li_110_450# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X95 hpd_0/negdff_0/ncsrl_0/a_n300_10# hpd_0/li_1860_2670# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X96 m1_n860_660# hpd_0/li_1860_2670# hpd_0/negdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.375 ps=3.5 w=0.5 l=0.5
X97 VSUBS hpd_0/negdff_0/li_110_450# hpd_0/negdff_0/m1_170_60# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X98 hpd_0/negdff_0/li_110_450# hpd_0/negdff_0/m1_170_60# hpd_0/negdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.5
X99 hpd_0/negdff_0/ncsrl_0/a_n470_450# m1_n8820_610# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X100 m1_n860_660# hpd_0/a_4100_2650# hpd_0/negdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X101 hpd_0/negdff_0/m1_170_60# m1_n8820_610# hpd_0/negdff_0/ncsrl_0/a_n300_n280# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X102 hpd_0/xor_0/a_n120_n150# hpd_0/li_3500_2650# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X103 hpd_0/xor_0/a_n120_n150# hpd_0/li_3500_2650# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X104 hpd_0/xor_0/a_n10_n310# hpd_0/a_4100_2650# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X105 hpd_0/xor_0/a_n10_n310# hpd_0/a_4100_2650# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X106 hpd_0/xor_0/a_n60_n280# hpd_0/xor_0/a_n120_n150# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.29625 ps=2.7 w=0.5 l=0.15
X107 m1_n920_n170# hpd_0/li_3500_2650# hpd_0/xor_0/a_n60_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29625 pd=2.7 as=0.1125 ps=0.95 w=0.5 l=0.15
X108 hpd_0/xor_0/a_n60_10# hpd_0/a_4100_2650# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.1125 pd=0.95 as=0.29625 ps=2.7 w=0.5 l=0.15
X109 m1_n920_n170# hpd_0/xor_0/a_n10_n310# hpd_0/xor_0/a_n60_n280# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29625 pd=2.7 as=0.0625 ps=0.75 w=0.5 l=0.15
X110 hpd_0/xor_0/a_n60_450# hpd_0/li_3500_2650# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1125 pd=0.95 as=0.29625 ps=2.7 w=0.5 l=0.15
X111 m1_n920_n170# hpd_0/xor_0/a_n10_n310# hpd_0/xor_0/a_n60_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.24625 pd=2.5 as=0.1125 ps=0.95 w=0.5 l=0.15
X112 hpd_0/xor_0/a_n60_740# hpd_0/a_4100_2650# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1125 pd=0.95 as=0.29625 ps=2.7 w=0.5 l=0.15
X113 m1_n920_n170# hpd_0/xor_0/a_n120_n150# hpd_0/xor_0/a_n60_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.24625 pd=2.5 as=0.1125 ps=0.95 w=0.5 l=0.15
X114 hpd_0/xor_1/a_n120_n150# hpd_0/a_460_2990# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X115 hpd_0/xor_1/a_n120_n150# hpd_0/a_460_2990# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X116 hpd_0/xor_1/a_n10_n310# hpd_0/a_4100_2650# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X117 hpd_0/xor_1/a_n10_n310# hpd_0/a_4100_2650# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X118 hpd_0/xor_1/a_n60_n280# hpd_0/xor_1/a_n120_n150# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.5 as=0 ps=0 w=0.5 l=0.15
X119 hpd_0/li_4860_2670# hpd_0/a_460_2990# hpd_0/xor_1/a_n60_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.5925 pd=5.4 as=0.225 ps=1.9 w=0.5 l=0.15
X120 hpd_0/xor_1/a_n60_10# hpd_0/a_4100_2650# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X121 hpd_0/li_4860_2670# hpd_0/xor_1/a_n10_n310# hpd_0/xor_1/a_n60_n280# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X122 hpd_0/xor_1/a_n60_450# hpd_0/a_460_2990# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0 ps=0 w=0.5 l=0.15
X123 hpd_0/li_4860_2670# hpd_0/xor_1/a_n10_n310# hpd_0/xor_1/a_n60_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.4925 pd=5 as=0 ps=0 w=0.5 l=0.15
X124 hpd_0/xor_1/a_n60_740# hpd_0/a_4100_2650# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.9 as=0 ps=0 w=0.5 l=0.15
X125 hpd_0/li_4860_2670# hpd_0/xor_1/a_n120_n150# hpd_0/xor_1/a_n60_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.15
X126 hpd_0/li_560_2670# hpd_0/a_460_2990# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X127 hpd_0/li_560_2670# hpd_0/a_460_2990# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X128 m1_n920_390# hpd_0/li_4860_2670# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X129 m1_n920_390# hpd_0/li_4860_2670# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X130 hpd_0/posdff_0/li_n550_450# hpd_0/posdff_0/m1_n490_60# hpd_0/posdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.375 ps=3.5 w=0.5 l=0.5
X131 hpd_0/posdff_0/csrl_0/a_n470_n150# m1_n8820_610# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.375 pd=3.5 as=0 ps=0 w=0.5 l=0.5
X132 hpd_0/posdff_0/csrl_0/a_n300_580# hpd_0/li_560_2670# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X133 hpd_0/posdff_0/csrl_0/a_n470_140# m1_n8820_610# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X134 m1_n860_660# hpd_0/posdff_0/m1_n490_60# hpd_0/posdff_0/li_n550_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X135 VSUBS hpd_0/a_460_2990# hpd_0/posdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X136 hpd_0/posdff_0/li_n550_450# m1_n8820_610# hpd_0/posdff_0/csrl_0/a_n300_580# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X137 hpd_0/posdff_0/csrl_0/a_n300_870# hpd_0/a_460_2990# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X138 hpd_0/posdff_0/m1_n490_60# hpd_0/posdff_0/li_n550_450# hpd_0/posdff_0/csrl_0/a_n470_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.5
X139 m1_n860_660# hpd_0/posdff_0/li_n550_450# hpd_0/posdff_0/m1_n490_60# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X140 VSUBS hpd_0/li_560_2670# hpd_0/posdff_0/csrl_0/a_n470_140# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X141 hpd_0/posdff_0/m1_n490_60# m1_n8820_610# hpd_0/posdff_0/csrl_0/a_n300_870# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X142 hpd_0/a_4100_2650# hpd_0/li_1860_2670# hpd_0/posdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.375 ps=3.5 w=0.5 l=0.5
X143 hpd_0/posdff_0/ncsrl_0/a_n470_740# m1_n8820_610# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X144 hpd_0/li_1860_2670# m1_n8820_610# hpd_0/posdff_0/ncsrl_0/a_n300_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.5
X145 hpd_0/posdff_0/ncsrl_0/a_n300_n280# hpd_0/posdff_0/m1_n490_60# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0 ps=0 w=0.5 l=0.5
X146 VSUBS hpd_0/a_4100_2650# hpd_0/li_1860_2670# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X147 hpd_0/posdff_0/ncsrl_0/a_n300_10# hpd_0/posdff_0/li_n550_450# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X148 m1_n860_660# hpd_0/posdff_0/li_n550_450# hpd_0/posdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.375 ps=3.5 w=0.5 l=0.5
X149 VSUBS hpd_0/li_1860_2670# hpd_0/a_4100_2650# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2 ps=1.8 w=0.5 l=0.5
X150 hpd_0/li_1860_2670# hpd_0/a_4100_2650# hpd_0/posdff_0/ncsrl_0/a_n470_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.5
X151 hpd_0/posdff_0/ncsrl_0/a_n470_450# m1_n8820_610# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X152 m1_n860_660# hpd_0/posdff_0/m1_n490_60# hpd_0/posdff_0/ncsrl_0/a_n470_740# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X153 hpd_0/a_4100_2650# m1_n8820_610# hpd_0/posdff_0/ncsrl_0/a_n300_n280# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X154 ipump_0/a_n180_450# li_n50_440# ipump_0/a_n260_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X155 ipump_0/a_n180_10# m1_n60_340# ipump_0/a_n260_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X156 m1_n150_240# m1_n920_n170# ipump_0/a_n20_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.15
X157 ipump_0/a_n340_450# li_n50_440# ipump_0/a_n420_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X158 ipump_0/a_n420_10# m1_n60_340# ipump_0/a_n500_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X159 ipump_0/a_n420_450# li_n50_440# ipump_0/a_n500_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X160 ipump_0/a_n20_450# li_n50_440# ipump_0/a_n100_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X161 ipump_0/a_n260_10# m1_n60_340# ipump_0/a_n340_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X162 ipump_0/a_n20_10# m1_n60_340# ipump_0/a_n100_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X163 m1_n150_240# m1_n920_390# ipump_0/a_n20_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.15
X164 ipump_0/a_n500_450# li_n50_440# ipump_0/a_n580_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X165 ipump_0/a_n500_10# m1_n60_340# ipump_0/a_n580_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X166 ipump_0/a_n100_10# m1_n60_340# ipump_0/a_n180_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X167 ipump_0/a_n100_450# li_n50_440# ipump_0/a_n180_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X168 ipump_0/a_n580_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.15
X169 ipump_0/a_n340_10# m1_n60_340# ipump_0/a_n420_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X170 ipump_0/a_n260_450# li_n50_440# ipump_0/a_n340_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.0625 pd=0.75 as=0.0625 ps=0.75 w=0.5 l=0.15
X171 ipump_0/a_n580_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.15
X172 vco_0/li_4880_260# vco_0/li_4480_260# vco_0/csi_11/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.15 ps=1.35 w=1 l=0.15
X173 vco_0/csi_11/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.35 as=0.175 ps=1.7 w=0.5 l=0.5
X174 vco_0/csi_11/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.35 as=0.175 ps=1.7 w=0.5 l=0.5
X175 vco_0/li_4880_260# vco_0/li_4480_260# vco_0/csi_11/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0.15 ps=1.35 w=1 l=0.15
X176 vco_0/li_4480_260# vco_0/li_4080_260# vco_0/csi_10/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X177 vco_0/csi_10/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X178 vco_0/csi_10/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X179 vco_0/li_4480_260# vco_0/li_4080_260# vco_0/csi_10/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X180 vco_0/li_130_240# vco_0/li_4880_260# vco_0/csi_12/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X181 vco_0/csi_12/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X182 vco_0/csi_12/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X183 vco_0/li_130_240# vco_0/li_4880_260# vco_0/csi_12/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X184 vco_0/li_480_260# vco_0/li_130_240# vco_0/csi_0/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X185 vco_0/csi_0/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X186 vco_0/csi_0/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X187 vco_0/li_480_260# vco_0/li_130_240# vco_0/csi_0/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X188 vco_0/li_880_260# vco_0/li_480_260# vco_0/csi_1/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X189 vco_0/csi_1/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X190 vco_0/csi_1/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X191 vco_0/li_880_260# vco_0/li_480_260# vco_0/csi_1/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X192 vco_0/li_1280_260# vco_0/li_880_260# vco_0/csi_2/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X193 vco_0/csi_2/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X194 vco_0/csi_2/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X195 vco_0/li_1280_260# vco_0/li_880_260# vco_0/csi_2/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X196 vco_0/li_2080_260# vco_0/li_1680_260# vco_0/csi_4/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X197 vco_0/csi_4/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X198 vco_0/csi_4/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X199 vco_0/li_2080_260# vco_0/li_1680_260# vco_0/csi_4/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X200 vco_0/li_1680_260# vco_0/li_1280_260# vco_0/csi_3/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X201 vco_0/csi_3/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X202 vco_0/csi_3/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X203 vco_0/li_1680_260# vco_0/li_1280_260# vco_0/csi_3/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X204 vco_0/li_2480_260# vco_0/li_2080_260# vco_0/csi_5/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X205 vco_0/csi_5/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X206 vco_0/csi_5/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X207 vco_0/li_2480_260# vco_0/li_2080_260# vco_0/csi_5/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X208 vco_0/li_2880_260# vco_0/li_2480_260# vco_0/csi_6/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X209 vco_0/csi_6/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X210 vco_0/csi_6/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X211 vco_0/li_2880_260# vco_0/li_2480_260# vco_0/csi_6/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X212 vco_0/li_3280_260# vco_0/li_2880_260# vco_0/csi_7/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X213 vco_0/csi_7/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X214 vco_0/csi_7/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X215 vco_0/li_3280_260# vco_0/li_2880_260# vco_0/csi_7/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X216 vco_0/li_3680_260# vco_0/li_3280_260# vco_0/csi_8/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X217 vco_0/csi_8/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X218 vco_0/csi_8/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X219 vco_0/li_3680_260# vco_0/li_3280_260# vco_0/csi_8/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X220 vco_0/li_4080_260# vco_0/li_3680_260# vco_0/csi_9/a_n40_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.7 as=0.3 ps=2.7 w=1 l=0.15
X221 vco_0/csi_9/a_n40_450# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=0.5 l=0.5
X222 vco_0/csi_9/a_n40_10# m1_n60_340# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X223 vco_0/li_4080_260# vco_0/li_3680_260# vco_0/csi_9/a_n40_450# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.7 as=0 ps=0 w=1 l=0.15
X224 vco_0/li_5510_260# vco_0/li_130_240# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X225 vco_0/li_5510_260# vco_0/li_130_240# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X226 m1_n9990_330# vco_0/li_5510_260# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X227 m1_n9990_330# vco_0/li_5510_260# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0 ps=0 w=0.5 l=0.15
X228 li_n50_440# m1_n150_240# vco_0/a_n1790_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.7 as=0.1 ps=0.9 w=0.5 l=0.5
X229 m1_n860_660# li_n50_440# li_n50_440# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.175 ps=1.7 w=0.5 l=0.5
X230 VSUBS m1_n60_340# m1_n60_340# VSUBS sky130_fd_pr__nfet_01v8 ad=0.025 pd=1.1 as=0.175 ps=1.7 w=0.5 l=0.5
X231 vco_0/a_n1790_10# m1_n150_240# li_n50_440# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X232 vco_0/a_n1790_10# m1_n150_240# li_n50_440# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X233 m1_n860_660# li_n50_440# li_n50_440# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X234 li_n50_440# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X235 li_n50_440# m1_n150_240# vco_0/a_n1790_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X236 li_n50_440# m1_n150_240# vco_0/a_n1790_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X237 m1_n860_660# li_n50_440# li_n50_440# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X238 li_n50_440# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X239 li_n50_440# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.175 pd=1.7 as=0.1 ps=0.9 w=0.5 l=0.5
X240 vco_0/a_n1790_10# m1_n150_240# li_n50_440# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X241 vco_0/a_n1790_10# m1_n150_240# li_n50_440# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X242 m1_n860_660# li_n50_440# li_n50_440# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X243 m1_n860_660# li_n50_440# m1_n60_340# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.025 pd=1.1 as=0.175 ps=1.7 w=0.5 l=0.5
X244 li_n50_440# m1_n150_240# vco_0/a_n1790_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X245 li_n50_440# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X246 li_n50_440# m1_n150_240# vco_0/a_n1790_10# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X247 m1_n860_660# li_n50_440# li_n50_440# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
X248 vco_0/a_n1790_10# m1_n150_240# li_n50_440# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.175 ps=1.7 w=0.5 l=0.5
X249 li_n50_440# li_n50_440# m1_n860_660# m1_n860_660# sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.5
C0 div8_0/div_2/li_100_660# m1_n860_660# 1.00934f
C1 m1_n860_660# m1_n8820_610# 3.85824f
C2 m1_n860_660# hpd_0/li_3500_2650# 1.22328f
C3 m1_n860_660# li_n50_440# 5.21046f
C4 vco_0/li_130_240# m1_n9990_330# 1.93015f
C5 m1_n150_240# li_n50_440# 1.04888f
C6 m1_n860_660# hpd_0/a_4100_2650# 1.30803f
C7 hpd_0/a_460_2990# m1_n860_660# 2.59074f
C8 VSUBS hpd_0/a_4100_2650# 1.04426f
C9 m1_n860_660# m1_n9990_330# 2.19963f
C10 m1_n60_340# 0 4.42575f **FLOATING
C11 li_n50_440# 0 3.48819f **FLOATING
C12 vco_0/li_130_240# 0 1.56669f **FLOATING
C13 m1_n150_240# 0 2.02737f **FLOATING
C14 hpd_0/a_4100_2650# 0 2.63709f **FLOATING
C15 m1_n8820_610# 0 4.7076f **FLOATING
C16 hpd_0/a_460_2990# 0 2.09549f **FLOATING
C17 hpd_0/negdff_0/m1_170_60# 0 1.08034f **FLOATING
C18 div8_0/div_2/li_100_660# 0 1.57707f **FLOATING
C19 div8_0/div_2/li_220_670# 0 1.27431f **FLOATING
C20 div8_0/m1_4560_860# 0 1.38577f **FLOATING
C21 div8_0/div_1/li_100_660# 0 1.57707f **FLOATING
C22 div8_0/div_1/li_220_670# 0 1.27431f **FLOATING
C23 m1_n860_660# 0 26.66077f **FLOATING
C24 div8_0/div_0/li_100_660# 0 1.57707f **FLOATING
C25 VSUBS 0 1.26832f **FLOATING
C26 div8_0/div_0/li_220_670# 0 1.27431f **FLOATING
C27 m1_n9990_330# 0 2.25355f **FLOATING
