magic
tech sky130A
timestamp 1765346561
<< nwell >>
rect -115 480 95 500
rect 85 420 95 440
<< locali >>
rect 55 225 135 245
<< metal1 >>
rect -115 480 95 500
rect 85 420 95 440
rect 55 225 135 245
rect 85 30 95 50
rect 65 -30 185 -10
use ext2spi  csrl_0
timestamp 1765332816
transform 1 0 330 0 1 30
box -255 -105 85 505
use ncsrl  ncsrl_0
timestamp 1765332714
transform 1 0 0 0 1 95
box -255 -155 85 450
<< end >>
