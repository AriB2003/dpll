magic
tech sky130A
timestamp 1765328216
<< nwell >>
rect -2845 540 -2665 640
rect 3735 545 3880 640
rect -4410 470 -2755 490
rect -4410 305 -4390 470
rect -2785 425 -2755 470
rect -535 330 -410 350
rect -480 220 -430 240
rect -25 220 10 240
rect -480 200 -460 220
<< locali >>
rect -2785 455 -2755 465
rect -2785 435 -2780 455
rect -2760 435 -2755 455
rect -2785 425 -2755 435
rect -535 330 -410 350
rect -535 315 -515 330
rect -430 315 -410 330
rect -480 220 -430 240
rect -25 220 10 240
rect -480 200 -460 220
rect -430 140 -390 145
rect -430 120 -420 140
rect -400 120 -390 140
rect -430 115 -390 120
rect -535 30 -515 45
rect -430 30 -410 45
rect -535 10 -410 30
<< viali >>
rect -2780 435 -2760 455
rect -420 120 -400 140
<< metal1 >>
rect -4410 470 -2755 490
rect -4410 305 -4390 470
rect -2785 455 -2755 470
rect -2785 435 -2780 455
rect -2760 435 -2755 455
rect -2785 425 -2755 435
rect -430 330 125 350
rect 95 315 125 330
rect -30 170 965 190
rect -430 140 -390 145
rect -430 120 -420 140
rect -400 120 -390 140
rect -75 120 50 140
rect -430 115 -390 120
rect -430 -65 -410 115
rect -385 10 1055 30
rect -460 -85 -410 -65
use div8  div8_0
timestamp 1765328216
transform 1 0 -5895 0 1 -260
box 700 20 3075 905
use hpd  hpd_0
timestamp 1765328216
transform 1 0 -3005 0 1 -1165
box 175 925 2565 1810
use ipump  ipump_0
timestamp 1765327476
transform 1 0 -90 0 1 40
box -360 -80 85 400
use vco  vco_0
timestamp 1765328216
transform 1 0 985 0 1 40
box -1000 -280 2895 605
<< end >>
