magic
tech sky130A
timestamp 1765330714
<< nwell >>
rect -360 140 85 300
<< nmos >>
rect -305 5 -290 55
rect -265 5 -250 55
rect -225 5 -210 55
rect -185 5 -170 55
rect -145 5 -130 55
rect -105 5 -90 55
rect -65 5 -50 55
rect -25 5 -10 55
rect 15 5 30 55
<< pmos >>
rect -305 225 -290 275
rect -265 225 -250 275
rect -225 225 -210 275
rect -185 225 -170 275
rect -145 225 -130 275
rect -105 225 -90 275
rect -65 225 -50 275
rect -25 225 -10 275
rect 15 225 30 275
<< ndiff >>
rect -340 40 -305 55
rect -340 20 -335 40
rect -315 20 -305 40
rect -340 5 -305 20
rect -290 5 -265 55
rect -250 5 -225 55
rect -210 5 -185 55
rect -170 5 -145 55
rect -130 5 -105 55
rect -90 5 -65 55
rect -50 5 -25 55
rect -10 5 15 55
rect 30 40 65 55
rect 30 20 40 40
rect 60 20 65 40
rect 30 5 65 20
<< pdiff >>
rect -340 260 -305 275
rect -340 240 -335 260
rect -315 240 -305 260
rect -340 225 -305 240
rect -290 225 -265 275
rect -250 225 -225 275
rect -210 225 -185 275
rect -170 225 -145 275
rect -130 225 -105 275
rect -90 225 -65 275
rect -50 225 -25 275
rect -10 225 15 275
rect 30 260 65 275
rect 30 240 40 260
rect 60 240 65 260
rect 30 225 65 240
<< ndiffc >>
rect -335 20 -315 40
rect 40 20 60 40
<< pdiffc >>
rect -335 240 -315 260
rect 40 240 60 260
<< psubdiff >>
rect -305 110 -255 115
rect -305 90 -290 110
rect -270 90 -255 110
rect -305 85 -255 90
<< nsubdiff >>
rect -305 190 -255 195
rect -305 170 -290 190
rect -270 170 -255 190
rect -305 165 -255 170
<< psubdiffcont >>
rect -290 90 -270 110
<< nsubdiffcont >>
rect -290 170 -270 190
<< poly >>
rect -305 285 -10 300
rect -305 275 -290 285
rect -265 275 -250 285
rect -225 275 -210 285
rect -185 275 -170 285
rect -145 275 -130 285
rect -105 275 -90 285
rect -65 275 -50 285
rect -25 275 -10 285
rect 15 275 30 290
rect -305 210 -290 225
rect -265 210 -250 225
rect -225 210 -210 225
rect -185 210 -170 225
rect -145 205 -130 225
rect -105 205 -90 225
rect -65 210 -50 225
rect -25 210 -10 225
rect -145 200 -90 205
rect -145 180 -120 200
rect -100 180 -90 200
rect -145 175 -90 180
rect -65 180 -25 185
rect 15 180 30 225
rect -65 160 -55 180
rect -35 165 30 180
rect -35 160 -25 165
rect -65 155 -25 160
rect -65 120 -25 125
rect -145 100 -90 105
rect -145 80 -120 100
rect -100 80 -90 100
rect -65 100 -55 120
rect -35 115 -25 120
rect -35 100 30 115
rect -65 95 -25 100
rect -145 75 -90 80
rect -305 55 -290 70
rect -265 55 -250 70
rect -225 55 -210 70
rect -185 55 -170 70
rect -145 55 -130 75
rect -105 55 -90 75
rect -65 55 -50 70
rect -25 55 -10 70
rect 15 55 30 100
rect -305 -5 -290 5
rect -265 -5 -250 5
rect -225 -5 -210 5
rect -185 -5 -170 5
rect -145 -5 -130 5
rect -105 -5 -90 5
rect -65 -5 -50 5
rect -25 -5 -10 5
rect -305 -20 -10 -5
rect 15 -10 30 5
<< polycont >>
rect -120 180 -100 200
rect -55 160 -35 180
rect -120 80 -100 100
rect -55 100 -35 120
<< locali >>
rect -340 260 -310 275
rect -340 240 -335 260
rect -315 240 -310 260
rect -340 225 -310 240
rect 35 260 65 270
rect 35 240 40 260
rect 60 240 65 260
rect 35 225 65 240
rect -330 195 -310 225
rect -130 205 15 225
rect -130 200 -90 205
rect -330 190 -260 195
rect -330 175 -290 190
rect -300 170 -290 175
rect -270 170 -260 190
rect -130 180 -120 200
rect -100 180 -90 200
rect -5 200 15 205
rect -130 175 -90 180
rect -65 180 -25 185
rect -5 180 65 200
rect -300 165 -260 170
rect -65 160 -55 180
rect -35 160 -25 180
rect -65 155 -25 160
rect 35 150 65 160
rect 35 130 40 150
rect 60 130 65 150
rect -65 120 -25 125
rect -300 110 -260 115
rect -300 90 -290 110
rect -270 90 -260 110
rect -300 85 -260 90
rect -130 100 -90 105
rect -290 55 -270 85
rect -130 80 -120 100
rect -100 80 -90 100
rect -65 100 -55 120
rect -35 100 -25 120
rect 35 100 65 130
rect -65 95 -25 100
rect -130 75 -90 80
rect -5 80 65 100
rect -5 75 15 80
rect -130 55 15 75
rect -340 40 -265 55
rect -340 20 -335 40
rect -315 20 -290 40
rect -270 20 -265 40
rect -340 5 -265 20
rect 35 40 65 55
rect 35 20 40 40
rect 60 20 65 40
rect 35 10 65 20
<< viali >>
rect -335 240 -315 260
rect 40 240 60 260
rect -55 160 -35 180
rect 40 130 60 150
rect -55 100 -35 120
rect -290 20 -270 40
rect 40 20 60 40
<< metal1 >>
rect -340 260 -310 300
rect -340 240 -335 260
rect -315 240 -310 260
rect -340 230 -310 240
rect -5 260 65 270
rect -5 240 40 260
rect 60 240 65 260
rect -5 225 65 240
rect -340 180 -25 185
rect -340 160 -55 180
rect -35 160 -25 180
rect -340 155 -25 160
rect -340 120 -25 125
rect -340 100 -55 120
rect -35 100 -25 120
rect -340 95 -25 100
rect -5 55 15 225
rect 35 150 65 160
rect 35 130 40 150
rect 60 130 65 150
rect 35 120 65 130
rect -295 40 -265 50
rect -295 20 -290 40
rect -270 20 -265 40
rect -295 -25 -265 20
rect -5 40 65 55
rect -5 20 40 40
rect 60 20 65 40
rect -5 10 65 20
<< end >>
