magic
tech sky130A
timestamp 1765304971
<< nwell >>
rect -145 530 35 605
rect -145 465 75 530
rect -295 140 85 465
<< nmos >>
rect -200 5 -150 55
rect -110 5 -60 55
rect -20 5 30 55
rect -200 -140 -150 -90
rect -110 -140 -60 -90
rect -20 -140 30 -90
<< pmos >>
rect -200 370 -150 420
rect -110 370 -60 420
rect -20 370 30 420
rect -200 225 -150 275
rect -110 225 -60 275
rect -20 225 30 275
<< ndiff >>
rect -235 5 -200 55
rect -150 5 -110 55
rect -60 40 -20 55
rect -60 20 -50 40
rect -30 20 -20 40
rect -60 5 -20 20
rect 30 5 65 55
rect -235 -90 -220 5
rect 50 -90 65 5
rect -235 -105 -200 -90
rect -235 -125 -230 -105
rect -210 -125 -200 -105
rect -235 -140 -200 -125
rect -150 -140 -110 -90
rect -60 -105 -20 -90
rect -60 -125 -50 -105
rect -30 -125 -20 -105
rect -60 -140 -20 -125
rect 30 -105 65 -90
rect 30 -125 40 -105
rect 60 -125 65 -105
rect 30 -140 65 -125
<< pdiff >>
rect -235 405 -200 420
rect -235 385 -230 405
rect -210 385 -200 405
rect -235 370 -200 385
rect -150 400 -110 420
rect -150 380 -140 400
rect -120 380 -110 400
rect -150 370 -110 380
rect -60 405 -20 420
rect -60 385 -50 405
rect -30 385 -20 405
rect -60 370 -20 385
rect 30 405 65 420
rect 30 385 40 405
rect 60 385 65 405
rect 30 370 65 385
rect -140 275 -120 370
rect -235 260 -200 275
rect -235 240 -230 260
rect -210 240 -200 260
rect -235 225 -200 240
rect -150 225 -110 275
rect -60 260 -20 275
rect -60 240 -50 260
rect -30 240 -20 260
rect -60 225 -20 240
rect 30 260 65 275
rect 30 240 40 260
rect 60 240 65 260
rect 30 225 65 240
<< ndiffc >>
rect -50 20 -30 40
rect -230 -125 -210 -105
rect -50 -125 -30 -105
rect 40 -125 60 -105
<< pdiffc >>
rect -230 385 -210 405
rect -140 380 -120 400
rect -50 385 -30 405
rect 40 385 60 405
rect -230 240 -210 260
rect -50 240 -30 260
rect 40 240 60 260
<< psubdiff >>
rect -20 -220 30 -205
rect -20 -245 -5 -220
rect 15 -245 30 -220
rect -20 -260 30 -245
<< nsubdiff >>
rect 5 495 55 510
rect 5 470 20 495
rect 40 470 55 495
rect 5 455 55 470
<< psubdiffcont >>
rect -5 -245 15 -220
<< nsubdiffcont >>
rect 20 470 40 495
<< poly >>
rect -200 420 -150 435
rect -110 420 -60 435
rect -20 420 30 435
rect -200 355 -150 370
rect -200 345 -170 355
rect -200 325 -195 345
rect -175 325 -170 345
rect -200 315 -170 325
rect -200 275 -150 290
rect -110 355 -60 370
rect -20 355 30 370
rect -95 290 -75 355
rect 15 345 65 355
rect 15 340 40 345
rect 35 325 40 340
rect 60 325 65 345
rect 35 315 65 325
rect -110 275 -60 290
rect -20 275 30 290
rect -200 210 -150 225
rect -110 210 -60 225
rect -20 210 30 225
rect -185 160 -165 210
rect -95 160 -75 210
rect -15 200 15 210
rect -15 180 -10 200
rect 10 180 15 200
rect -15 170 15 180
rect -195 150 -165 160
rect -195 130 -190 150
rect -170 130 -165 150
rect -195 120 -165 130
rect -105 150 -75 160
rect -105 130 -100 150
rect -80 130 -75 150
rect -105 120 -75 130
rect -185 70 -165 120
rect -95 70 -75 120
rect -15 100 15 110
rect -15 80 -10 100
rect 10 80 15 100
rect -15 70 15 80
rect -200 55 -150 70
rect -110 55 -60 70
rect -20 55 30 70
rect -200 -10 -150 5
rect -110 -10 -60 5
rect -20 -10 30 5
rect -200 -45 -170 -35
rect -200 -65 -195 -45
rect -175 -65 -170 -45
rect -200 -75 -170 -65
rect -95 -75 -75 -10
rect 0 -45 30 -35
rect 0 -65 5 -45
rect 25 -65 30 -45
rect 0 -75 30 -65
rect -200 -90 -150 -75
rect -110 -90 -60 -75
rect -20 -90 30 -75
rect -200 -155 -150 -140
rect -110 -155 -60 -140
rect -20 -155 30 -140
<< polycont >>
rect -195 325 -175 345
rect 40 325 60 345
rect -10 180 10 200
rect -190 130 -170 150
rect -100 130 -80 150
rect -10 80 10 100
rect -195 -65 -175 -45
rect 5 -65 25 -45
<< locali >>
rect 15 495 45 505
rect 15 470 20 495
rect 40 470 45 495
rect 15 460 45 470
rect -225 430 -35 450
rect -225 415 -205 430
rect -235 405 -205 415
rect -55 415 -35 430
rect -235 385 -230 405
rect -210 385 -205 405
rect -235 375 -205 385
rect -145 400 -115 410
rect -145 380 -140 400
rect -120 380 -115 400
rect -145 370 -115 380
rect -55 405 -25 415
rect -55 385 -50 405
rect -30 385 -25 405
rect 35 405 65 415
rect 35 395 40 405
rect -55 375 -25 385
rect -5 385 40 395
rect 60 385 65 405
rect -5 375 65 385
rect -200 345 -170 355
rect -200 325 -195 345
rect -175 325 -170 345
rect -200 315 -170 325
rect -235 260 -205 270
rect -235 240 -230 260
rect -210 250 -205 260
rect -55 260 -25 270
rect -55 250 -50 260
rect -210 240 -50 250
rect -30 240 -25 260
rect -235 230 -25 240
rect -5 210 15 375
rect -15 200 15 210
rect -15 180 -10 200
rect 10 180 15 200
rect -15 170 15 180
rect -195 150 -165 160
rect -235 130 -190 150
rect -170 130 -165 150
rect -195 120 -165 130
rect -105 150 -75 160
rect -105 130 -100 150
rect -80 130 -75 150
rect -105 120 -75 130
rect -5 110 15 170
rect -15 100 15 110
rect -15 90 -10 100
rect -95 80 -10 90
rect 10 80 15 100
rect -95 70 15 80
rect 35 345 65 355
rect 35 325 40 345
rect 60 325 65 345
rect 35 315 65 325
rect 35 270 55 315
rect 35 260 65 270
rect 35 240 40 260
rect 60 240 65 260
rect 35 230 65 240
rect 35 150 55 230
rect 35 130 85 150
rect -95 -10 -75 70
rect -55 40 -25 50
rect -55 20 -50 40
rect -30 30 -25 40
rect 35 30 55 130
rect -30 20 55 30
rect -55 10 55 20
rect -95 -30 -35 -10
rect -200 -45 -170 -35
rect -200 -65 -195 -45
rect -175 -65 -170 -45
rect -200 -75 -170 -65
rect -55 -95 -35 -30
rect 0 -35 20 10
rect 0 -45 30 -35
rect 0 -65 5 -45
rect 25 -65 30 -45
rect 0 -75 30 -65
rect -235 -105 -205 -95
rect -235 -125 -230 -105
rect -210 -125 -205 -105
rect -235 -135 -205 -125
rect -55 -105 -25 -95
rect -55 -125 -50 -105
rect -30 -125 -25 -105
rect -55 -140 -25 -125
rect 35 -105 65 -95
rect 35 -125 40 -105
rect 60 -125 65 -105
rect 35 -135 65 -125
rect -10 -220 20 -210
rect -10 -245 -5 -220
rect 15 -245 20 -220
rect -10 -255 20 -245
<< viali >>
rect -140 380 -120 400
rect -195 325 -175 345
rect -10 180 10 200
rect -100 130 -80 150
rect -10 80 10 100
rect -195 -65 -175 -45
rect -230 -125 -210 -105
rect 40 -125 60 -105
<< metal1 >>
rect -145 400 -115 410
rect -145 380 -140 400
rect -120 380 -115 400
rect -145 370 -115 380
rect -200 345 -170 355
rect -235 325 -195 345
rect -175 325 -170 345
rect -200 315 -170 325
rect -5 325 85 345
rect -5 210 15 325
rect -15 200 15 210
rect -15 180 -10 200
rect 10 180 15 200
rect -15 170 15 180
rect -105 150 -75 160
rect -235 130 -100 150
rect -80 130 85 150
rect -105 120 -75 130
rect -15 100 15 110
rect -15 80 -10 100
rect 10 80 15 100
rect -15 70 15 80
rect -200 -45 -170 -35
rect -235 -65 -195 -45
rect -175 -65 -170 -45
rect -5 -45 15 70
rect -5 -65 85 -45
rect -200 -75 -170 -65
rect -235 -105 -205 -95
rect 35 -105 65 -95
rect -235 -125 -230 -105
rect -210 -125 40 -105
rect 60 -125 65 -105
rect -235 -135 -205 -125
rect 35 -135 65 -125
<< end >>
