magic
tech sky130A
timestamp 1765307270
<< nwell >>
rect -295 205 85 640
<< nmos >>
rect -200 70 -150 120
rect -110 70 -60 120
rect -20 70 30 120
rect -200 -75 -150 -25
rect -110 -75 -60 -25
rect -20 -75 30 -25
<< pmos >>
rect -200 435 -150 485
rect -110 435 -60 485
rect -20 435 30 485
rect -200 290 -150 340
rect -110 290 -60 340
rect -20 290 30 340
<< ndiff >>
rect -235 105 -200 120
rect -235 85 -230 105
rect -210 85 -200 105
rect -235 70 -200 85
rect -150 70 -110 120
rect -60 105 -20 120
rect -60 85 -50 105
rect -30 85 -20 105
rect -60 70 -20 85
rect 30 105 65 120
rect 30 85 40 105
rect 60 85 65 105
rect 30 70 65 85
rect -140 -25 -120 70
rect -235 -40 -200 -25
rect -235 -60 -230 -40
rect -210 -60 -200 -40
rect -235 -75 -200 -60
rect -150 -35 -110 -25
rect -150 -55 -140 -35
rect -120 -55 -110 -35
rect -150 -75 -110 -55
rect -60 -40 -20 -25
rect -60 -60 -50 -40
rect -30 -60 -20 -40
rect -60 -75 -20 -60
rect 30 -40 65 -25
rect 30 -60 40 -40
rect 60 -60 65 -40
rect 30 -75 65 -60
<< pdiff >>
rect -235 470 -200 485
rect -235 450 -230 470
rect -210 450 -200 470
rect -235 435 -200 450
rect -150 435 -110 485
rect -60 470 -20 485
rect -60 450 -50 470
rect -30 450 -20 470
rect -60 435 -20 450
rect 30 470 65 485
rect 30 450 40 470
rect 60 450 65 470
rect 30 435 65 450
rect -235 340 -220 435
rect 50 340 65 435
rect -235 290 -200 340
rect -150 290 -110 340
rect -60 325 -20 340
rect -60 305 -50 325
rect -30 305 -20 325
rect -60 290 -20 305
rect 30 290 65 340
<< ndiffc >>
rect -230 85 -210 105
rect -50 85 -30 105
rect 40 85 60 105
rect -230 -60 -210 -40
rect -140 -55 -120 -35
rect -50 -60 -30 -40
rect 40 -60 60 -40
<< pdiffc >>
rect -230 450 -210 470
rect -50 450 -30 470
rect 40 450 60 470
rect -50 305 -30 325
<< psubdiff >>
rect 5 -125 55 -110
rect 5 -150 20 -125
rect 40 -150 55 -125
rect 5 -165 55 -150
<< nsubdiff >>
rect -20 590 30 605
rect -20 565 -5 590
rect 15 565 30 590
rect -20 550 30 565
<< psubdiffcont >>
rect 20 -150 40 -125
<< nsubdiffcont >>
rect -5 565 15 590
<< poly >>
rect -200 485 -150 500
rect -110 485 -60 500
rect -20 485 30 500
rect -200 420 -150 435
rect -110 420 -60 435
rect -20 420 30 435
rect -200 410 -170 420
rect -200 390 -195 410
rect -175 390 -170 410
rect -200 380 -170 390
rect -95 355 -75 420
rect 0 410 30 420
rect 0 390 5 410
rect 25 390 30 410
rect 0 380 30 390
rect -200 340 -150 355
rect -110 340 -60 355
rect -20 340 30 355
rect -200 275 -150 290
rect -110 275 -60 290
rect -20 275 30 290
rect -185 225 -165 275
rect -95 225 -75 275
rect -15 265 15 275
rect -15 245 -10 265
rect 10 245 15 265
rect -15 235 15 245
rect -195 215 -165 225
rect -195 195 -190 215
rect -170 195 -165 215
rect -195 185 -165 195
rect -105 215 -75 225
rect -105 195 -100 215
rect -80 195 -75 215
rect -105 185 -75 195
rect -185 135 -165 185
rect -95 135 -75 185
rect -15 165 15 175
rect -15 145 -10 165
rect 10 145 15 165
rect -15 135 15 145
rect -200 120 -150 135
rect -110 120 -60 135
rect -20 120 30 135
rect -200 55 -150 70
rect -200 20 -170 30
rect -200 0 -195 20
rect -175 0 -170 20
rect -200 -10 -170 0
rect -200 -25 -150 -10
rect -110 55 -60 70
rect -20 55 30 70
rect -95 -10 -75 55
rect 35 20 65 30
rect 35 5 40 20
rect 15 0 40 5
rect 60 0 65 20
rect 15 -10 65 0
rect -110 -25 -60 -10
rect -20 -25 30 -10
rect -200 -90 -150 -75
rect -110 -90 -60 -75
rect -20 -90 30 -75
<< polycont >>
rect -195 390 -175 410
rect 5 390 25 410
rect -10 245 10 265
rect -190 195 -170 215
rect -100 195 -80 215
rect -10 145 10 165
rect -195 0 -175 20
rect 40 0 60 20
<< locali >>
rect -10 590 20 600
rect -10 565 -5 590
rect 15 565 20 590
rect -10 555 20 565
rect -235 470 -205 480
rect -235 450 -230 470
rect -210 450 -205 470
rect -235 440 -205 450
rect -55 470 -25 485
rect -55 450 -50 470
rect -30 450 -25 470
rect -55 440 -25 450
rect 35 470 65 480
rect 35 450 40 470
rect 60 450 65 470
rect 35 440 65 450
rect -200 410 -170 420
rect -200 390 -195 410
rect -175 390 -170 410
rect -200 380 -170 390
rect -55 375 -35 440
rect -95 355 -35 375
rect 0 410 30 420
rect 0 390 5 410
rect 25 390 30 410
rect 0 380 30 390
rect -95 275 -75 355
rect 0 335 20 380
rect -55 325 55 335
rect -55 305 -50 325
rect -30 315 55 325
rect -30 305 -25 315
rect -55 295 -25 305
rect -95 265 15 275
rect -95 255 -10 265
rect -15 245 -10 255
rect 10 245 15 265
rect -15 235 15 245
rect -195 215 -165 225
rect -195 195 -190 215
rect -170 195 -165 215
rect -195 185 -165 195
rect -105 215 -75 225
rect -105 195 -100 215
rect -80 195 -75 215
rect -105 185 -75 195
rect -5 175 15 235
rect -15 165 15 175
rect -15 145 -10 165
rect 10 145 15 165
rect -15 135 15 145
rect -235 105 -25 115
rect -235 85 -230 105
rect -210 95 -50 105
rect -210 85 -205 95
rect -235 75 -205 85
rect -55 85 -50 95
rect -30 85 -25 105
rect -55 75 -25 85
rect -200 20 -170 30
rect -200 0 -195 20
rect -175 0 -170 20
rect -200 -10 -170 0
rect -235 -40 -205 -30
rect -235 -60 -230 -40
rect -210 -60 -205 -40
rect -235 -70 -205 -60
rect -145 -35 -115 -25
rect -5 -30 15 135
rect 35 115 55 315
rect 35 105 65 115
rect 35 85 40 105
rect 60 85 65 105
rect 35 75 65 85
rect 35 30 55 75
rect 35 20 65 30
rect 35 0 40 20
rect 60 0 65 20
rect 35 -10 65 0
rect -145 -55 -140 -35
rect -120 -55 -115 -35
rect -145 -65 -115 -55
rect -55 -40 -25 -30
rect -55 -60 -50 -40
rect -30 -60 -25 -40
rect -5 -40 65 -30
rect -5 -50 40 -40
rect -225 -85 -205 -70
rect -55 -70 -25 -60
rect 35 -60 40 -50
rect 60 -60 65 -40
rect 35 -70 65 -60
rect -55 -85 -35 -70
rect -225 -105 -35 -85
rect 15 -125 45 -115
rect 15 -150 20 -125
rect 40 -150 45 -125
rect 15 -160 45 -150
<< viali >>
rect -230 450 -210 470
rect 40 450 60 470
rect -195 390 -175 410
rect -10 245 10 265
rect -100 195 -80 215
rect -10 145 10 165
rect -195 0 -175 20
rect -140 -55 -120 -35
<< metal1 >>
rect -235 470 -205 480
rect 35 470 65 480
rect -235 450 -230 470
rect -210 450 40 470
rect 60 450 65 470
rect -235 440 -205 450
rect 35 440 65 450
rect -200 410 -170 420
rect -235 390 -195 410
rect -175 390 -170 410
rect -200 380 -170 390
rect -5 390 85 410
rect -5 275 15 390
rect -15 265 15 275
rect -15 245 -10 265
rect 10 245 15 265
rect -15 235 15 245
rect -105 215 -75 225
rect -195 195 -100 215
rect -80 195 55 215
rect -105 185 -75 195
rect -15 165 15 175
rect -15 145 -10 165
rect 10 145 15 165
rect -15 135 15 145
rect -200 20 -170 30
rect -235 0 -195 20
rect -175 0 -170 20
rect -5 20 15 135
rect -5 0 85 20
rect -200 -10 -170 0
rect -145 -35 -115 -25
rect -145 -55 -140 -35
rect -120 -55 -115 -35
rect -145 -65 -115 -55
<< end >>
