magic
tech sky130A
timestamp 1765148092
<< nwell >>
rect -25 220 10 240
<< locali >>
rect -25 220 10 240
<< metal1 >>
rect -30 170 965 190
rect -75 120 50 140
use ipump  ipump_0
timestamp 1765147879
transform 1 0 -90 0 1 40
box -360 -80 85 400
use vco  vco_0
timestamp 1765143928
transform 1 0 985 0 1 40
box -1000 -85 2895 455
<< end >>
