magic
tech sky130A
magscale 1 2
timestamp 1765240007
<< error_p >>
rect -186 150 -180 166
rect -120 160 -60 170
rect -120 150 -114 160
rect -82 144 -60 160
rect -144 140 -120 144
rect -82 140 -30 144
rect -170 134 -154 140
rect -146 134 -130 140
rect -110 106 -50 110
rect -150 10 -96 34
rect -180 -35 -150 -20
<< nwell >>
rect -290 1060 70 1210
rect -290 930 150 1060
rect -290 280 170 930
<< nmos >>
rect -400 10 -300 110
rect -220 10 -120 110
rect -40 10 60 110
rect -400 -280 -300 -180
rect -220 -280 -120 -180
rect -40 -280 60 -180
<< pmos >>
rect -90 740 -60 840
rect 30 740 60 840
rect -90 450 -60 550
rect 30 450 60 550
<< ndiff >>
rect -470 80 -400 110
rect -470 40 -460 80
rect -420 40 -400 80
rect -470 10 -400 40
rect -300 80 -220 110
rect -300 40 -280 80
rect -240 40 -220 80
rect -300 10 -220 40
rect -120 80 -40 110
rect -120 40 -100 80
rect -60 40 -40 80
rect -120 10 -40 40
rect 60 80 130 110
rect 60 40 80 80
rect 120 40 130 80
rect 60 10 130 40
rect -470 -20 -440 10
rect -180 -50 -150 -20
rect -470 -180 -440 -150
rect 100 -180 130 10
rect -470 -210 -400 -180
rect -470 -250 -460 -210
rect -420 -250 -400 -210
rect -470 -280 -400 -250
rect -300 -210 -220 -180
rect -300 -250 -280 -210
rect -240 -250 -220 -210
rect -300 -280 -220 -250
rect -120 -210 -40 -180
rect -120 -250 -100 -210
rect -60 -250 -40 -210
rect -120 -280 -40 -250
rect 60 -210 130 -180
rect 60 -250 80 -210
rect 120 -250 130 -210
rect 60 -280 130 -250
<< pdiff >>
rect -180 810 -90 840
rect -180 770 -170 810
rect -130 770 -90 810
rect -180 740 -90 770
rect -60 740 30 840
rect 60 740 130 840
rect -180 550 -150 740
rect 100 550 130 740
rect -180 450 -90 550
rect -60 450 30 550
rect 60 520 130 550
rect 60 480 80 520
rect 120 480 130 520
rect 60 450 130 480
<< ndiffc >>
rect -460 40 -420 80
rect -280 40 -240 80
rect -100 40 -60 80
rect 80 40 120 80
rect -460 -250 -420 -210
rect -280 -250 -240 -210
rect -100 -250 -60 -210
rect 80 -250 120 -210
<< pdiffc >>
rect -170 770 -130 810
rect 80 480 120 520
<< psubdiff >>
rect -40 -440 60 -410
rect -40 -490 -10 -440
rect 30 -490 60 -440
rect -40 -520 60 -490
<< nsubdiff >>
rect 10 990 110 1020
rect 10 940 40 990
rect 80 940 110 990
rect 10 910 110 940
<< psubdiffcont >>
rect -10 -490 30 -440
<< nsubdiffcont >>
rect 40 940 80 990
<< poly >>
rect -90 840 -60 870
rect 30 840 60 870
rect -90 710 -60 740
rect 30 710 60 740
rect -90 550 -60 580
rect 30 550 60 580
rect -90 400 -60 450
rect 30 420 60 450
rect -180 370 -60 400
rect -90 280 -60 370
rect -10 400 60 420
rect -10 360 0 400
rect 40 360 60 400
rect -10 340 60 360
rect -90 250 60 280
rect -180 190 -120 210
rect -180 150 -170 190
rect -130 160 -120 190
rect -130 150 -60 160
rect -180 140 -60 150
rect 30 140 60 250
rect -400 110 -300 140
rect -220 110 -120 140
rect -40 110 60 140
rect -400 -20 -300 10
rect -220 -20 -120 10
rect -40 -20 60 10
rect -400 -180 -300 -150
rect -220 -180 -120 -150
rect -40 -180 60 -150
rect -400 -310 -300 -280
rect -220 -310 -120 -280
rect -40 -310 60 -280
<< polycont >>
rect 0 360 40 400
rect -170 150 -130 190
<< locali >>
rect 30 990 90 1010
rect 30 940 40 990
rect 80 940 90 990
rect 30 920 90 940
rect -180 810 -120 840
rect -180 770 -170 810
rect -130 770 -120 810
rect -180 750 -120 770
rect -170 210 -130 550
rect -10 500 30 550
rect -90 460 30 500
rect 70 520 130 550
rect 70 480 80 520
rect 120 480 130 520
rect -90 300 -50 460
rect 70 450 130 480
rect -10 400 50 420
rect -10 360 0 400
rect 40 360 50 400
rect -10 340 50 360
rect -90 260 -30 300
rect -180 190 -120 210
rect -180 150 -170 190
rect -130 150 -120 190
rect -180 140 -120 150
rect -70 140 -30 260
rect 10 140 50 340
rect -470 80 -410 110
rect -470 40 -460 80
rect -420 40 -410 80
rect -470 20 -410 40
rect -290 80 -230 110
rect -290 40 -280 80
rect -240 40 -230 80
rect -290 20 -230 40
rect -110 80 -50 110
rect -110 40 -100 80
rect -60 40 -50 80
rect -110 20 -50 40
rect 70 80 130 110
rect 70 40 80 80
rect 120 40 130 80
rect 70 20 130 40
rect -470 -210 -410 -190
rect -470 -250 -460 -210
rect -420 -250 -410 -210
rect -470 -280 -410 -250
rect -290 -210 -230 -190
rect -290 -250 -280 -210
rect -240 -250 -230 -210
rect -290 -280 -230 -250
rect -110 -210 -50 -190
rect -110 -250 -100 -210
rect -60 -250 -50 -210
rect -110 -280 -50 -250
rect 70 -210 130 -190
rect 70 -250 80 -210
rect 120 -250 130 -210
rect 70 -280 130 -250
rect -20 -440 40 -420
rect -20 -490 -10 -440
rect 30 -490 40 -440
rect -20 -510 40 -490
<< end >>
